-- system_disp_7_seg.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_disp_7_seg is
	port (
		pio_disp_0_clk_clk                    : in  std_logic                     := '0';             --                 pio_disp_0_clk.clk
		pio_disp_0_external_connection_export : out std_logic_vector(7 downto 0);                     -- pio_disp_0_external_connection.export
		pio_disp_0_reset_reset_n              : in  std_logic                     := '0';             --               pio_disp_0_reset.reset_n
		pio_disp_0_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  pio_disp_0_s1.address
		pio_disp_0_s1_write_n                 : in  std_logic                     := '0';             --                               .write_n
		pio_disp_0_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		pio_disp_0_s1_chipselect              : in  std_logic                     := '0';             --                               .chipselect
		pio_disp_0_s1_readdata                : out std_logic_vector(31 downto 0);                    --                               .readdata
		pio_disp_1_clk_clk                    : in  std_logic                     := '0';             --                 pio_disp_1_clk.clk
		pio_disp_1_external_connection_export : out std_logic_vector(7 downto 0);                     -- pio_disp_1_external_connection.export
		pio_disp_1_reset_reset_n              : in  std_logic                     := '0';             --               pio_disp_1_reset.reset_n
		pio_disp_1_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  pio_disp_1_s1.address
		pio_disp_1_s1_write_n                 : in  std_logic                     := '0';             --                               .write_n
		pio_disp_1_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		pio_disp_1_s1_chipselect              : in  std_logic                     := '0';             --                               .chipselect
		pio_disp_1_s1_readdata                : out std_logic_vector(31 downto 0);                    --                               .readdata
		pio_disp_2_clk_clk                    : in  std_logic                     := '0';             --                 pio_disp_2_clk.clk
		pio_disp_2_external_connection_export : out std_logic_vector(7 downto 0);                     -- pio_disp_2_external_connection.export
		pio_disp_2_reset_reset_n              : in  std_logic                     := '0';             --               pio_disp_2_reset.reset_n
		pio_disp_2_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  pio_disp_2_s1.address
		pio_disp_2_s1_write_n                 : in  std_logic                     := '0';             --                               .write_n
		pio_disp_2_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		pio_disp_2_s1_chipselect              : in  std_logic                     := '0';             --                               .chipselect
		pio_disp_2_s1_readdata                : out std_logic_vector(31 downto 0);                    --                               .readdata
		pio_disp_3_clk_clk                    : in  std_logic                     := '0';             --                 pio_disp_3_clk.clk
		pio_disp_3_external_connection_export : out std_logic_vector(7 downto 0);                     -- pio_disp_3_external_connection.export
		pio_disp_3_reset_reset_n              : in  std_logic                     := '0';             --               pio_disp_3_reset.reset_n
		pio_disp_3_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  pio_disp_3_s1.address
		pio_disp_3_s1_write_n                 : in  std_logic                     := '0';             --                               .write_n
		pio_disp_3_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		pio_disp_3_s1_chipselect              : in  std_logic                     := '0';             --                               .chipselect
		pio_disp_3_s1_readdata                : out std_logic_vector(31 downto 0);                    --                               .readdata
		pio_disp_4_clk_clk                    : in  std_logic                     := '0';             --                 pio_disp_4_clk.clk
		pio_disp_4_external_connection_export : out std_logic_vector(7 downto 0);                     -- pio_disp_4_external_connection.export
		pio_disp_4_reset_reset_n              : in  std_logic                     := '0';             --               pio_disp_4_reset.reset_n
		pio_disp_4_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  pio_disp_4_s1.address
		pio_disp_4_s1_write_n                 : in  std_logic                     := '0';             --                               .write_n
		pio_disp_4_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		pio_disp_4_s1_chipselect              : in  std_logic                     := '0';             --                               .chipselect
		pio_disp_4_s1_readdata                : out std_logic_vector(31 downto 0);                    --                               .readdata
		pio_disp_5_clk_clk                    : in  std_logic                     := '0';             --                 pio_disp_5_clk.clk
		pio_disp_5_external_connection_export : out std_logic_vector(7 downto 0);                     -- pio_disp_5_external_connection.export
		pio_disp_5_reset_reset_n              : in  std_logic                     := '0';             --               pio_disp_5_reset.reset_n
		pio_disp_5_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  pio_disp_5_s1.address
		pio_disp_5_s1_write_n                 : in  std_logic                     := '0';             --                               .write_n
		pio_disp_5_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		pio_disp_5_s1_chipselect              : in  std_logic                     := '0';             --                               .chipselect
		pio_disp_5_s1_readdata                : out std_logic_vector(31 downto 0)                     --                               .readdata
	);
end entity system_disp_7_seg;

architecture rtl of system_disp_7_seg is
	component system_disp_7_seg_pio_disp_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component system_disp_7_seg_pio_disp_0;

begin

	pio_disp_0 : component system_disp_7_seg_pio_disp_0
		port map (
			clk        => pio_disp_0_clk_clk,                    --                 clk.clk
			reset_n    => pio_disp_0_reset_reset_n,              --               reset.reset_n
			address    => pio_disp_0_s1_address,                 --                  s1.address
			write_n    => pio_disp_0_s1_write_n,                 --                    .write_n
			writedata  => pio_disp_0_s1_writedata,               --                    .writedata
			chipselect => pio_disp_0_s1_chipselect,              --                    .chipselect
			readdata   => pio_disp_0_s1_readdata,                --                    .readdata
			out_port   => pio_disp_0_external_connection_export  -- external_connection.export
		);

	pio_disp_1 : component system_disp_7_seg_pio_disp_0
		port map (
			clk        => pio_disp_1_clk_clk,                    --                 clk.clk
			reset_n    => pio_disp_1_reset_reset_n,              --               reset.reset_n
			address    => pio_disp_1_s1_address,                 --                  s1.address
			write_n    => pio_disp_1_s1_write_n,                 --                    .write_n
			writedata  => pio_disp_1_s1_writedata,               --                    .writedata
			chipselect => pio_disp_1_s1_chipselect,              --                    .chipselect
			readdata   => pio_disp_1_s1_readdata,                --                    .readdata
			out_port   => pio_disp_1_external_connection_export  -- external_connection.export
		);

	pio_disp_2 : component system_disp_7_seg_pio_disp_0
		port map (
			clk        => pio_disp_2_clk_clk,                    --                 clk.clk
			reset_n    => pio_disp_2_reset_reset_n,              --               reset.reset_n
			address    => pio_disp_2_s1_address,                 --                  s1.address
			write_n    => pio_disp_2_s1_write_n,                 --                    .write_n
			writedata  => pio_disp_2_s1_writedata,               --                    .writedata
			chipselect => pio_disp_2_s1_chipselect,              --                    .chipselect
			readdata   => pio_disp_2_s1_readdata,                --                    .readdata
			out_port   => pio_disp_2_external_connection_export  -- external_connection.export
		);

	pio_disp_3 : component system_disp_7_seg_pio_disp_0
		port map (
			clk        => pio_disp_3_clk_clk,                    --                 clk.clk
			reset_n    => pio_disp_3_reset_reset_n,              --               reset.reset_n
			address    => pio_disp_3_s1_address,                 --                  s1.address
			write_n    => pio_disp_3_s1_write_n,                 --                    .write_n
			writedata  => pio_disp_3_s1_writedata,               --                    .writedata
			chipselect => pio_disp_3_s1_chipselect,              --                    .chipselect
			readdata   => pio_disp_3_s1_readdata,                --                    .readdata
			out_port   => pio_disp_3_external_connection_export  -- external_connection.export
		);

	pio_disp_4 : component system_disp_7_seg_pio_disp_0
		port map (
			clk        => pio_disp_4_clk_clk,                    --                 clk.clk
			reset_n    => pio_disp_4_reset_reset_n,              --               reset.reset_n
			address    => pio_disp_4_s1_address,                 --                  s1.address
			write_n    => pio_disp_4_s1_write_n,                 --                    .write_n
			writedata  => pio_disp_4_s1_writedata,               --                    .writedata
			chipselect => pio_disp_4_s1_chipselect,              --                    .chipselect
			readdata   => pio_disp_4_s1_readdata,                --                    .readdata
			out_port   => pio_disp_4_external_connection_export  -- external_connection.export
		);

	pio_disp_5 : component system_disp_7_seg_pio_disp_0
		port map (
			clk        => pio_disp_5_clk_clk,                    --                 clk.clk
			reset_n    => pio_disp_5_reset_reset_n,              --               reset.reset_n
			address    => pio_disp_5_s1_address,                 --                  s1.address
			write_n    => pio_disp_5_s1_write_n,                 --                    .write_n
			writedata  => pio_disp_5_s1_writedata,               --                    .writedata
			chipselect => pio_disp_5_s1_chipselect,              --                    .chipselect
			readdata   => pio_disp_5_s1_readdata,                --                    .readdata
			out_port   => pio_disp_5_external_connection_export  -- external_connection.export
		);

end architecture rtl; -- of system_disp_7_seg
