00009197
80018193
00010117
ff810113
088000ef
0000006f
00000000
00000000
fe010113
00112e23
00812c23
00912a23
02010413
fea42623
fec42783
00078863
fec42703
00100793
00f71663
00100793
0300006f
fec42783
fff78793
00078513
fc1ff0ef
00050493
fec42783
ffe78793
00078513
fadff0ef
00050793
00f487b3
00078513
01c12083
01812403
01412483
02010113
00008067
fe010113
00112e23
00812c23
02010413
fe042623
0340006f
fec42503
f6dff0ef
00050693
000087b7
00078713
fec42783
00279793
00f707b3
00d7a023
fec42783
00178793
fef42623
fec42703
00900793
fce7d4e3
00000793
00078513
01c12083
01812403
02010113
00008067
