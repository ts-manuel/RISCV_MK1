00001197
80018193
20000517
42050513
20000617
47860613
40a60633
00000593
228000ef
00000517
47450513
00050863
00000517
41450513
460000ef
180000ef
00012503
00410593
00000613
0d4000ef
13c0006f
ff010113
00812423
20000437
44044783
00112623
02079263
00000793
00078a63
20000537
42850513
00000097
000000e7
00100793
44f40023
00c12083
00812403
01010113
00008067
00000793
00078e63
200005b7
20000537
44458593
42850513
00000317
00000067
00008067
fe010113
00112e23
00812c23
02010413
fea42623
fec42783
00078863
fec42703
00100793
00f71663
00100793
0200006f
fec42783
fff78793
00078513
fc5ff0ef
00050713
fec42783
00f707b3
00078513
01c12083
01812403
02010113
00008067
fe010113
00112e23
00812c23
02010413
fe042623
0340006f
fec42503
f85ff0ef
00050693
200007b7
45c78713
fec42783
00279793
00f707b3
00d7a023
fec42783
00178793
fef42623
fec42703
00900793
fce7d4e3
00000793
00078513
01c12083
01812403
02010113
00008067
ff010113
00000593
00812423
00112623
00050413
184000ef
59402503
03c52783
00078463
000780e7
00040513
38c000ef
ff010113
00812423
01212023
00000793
00000913
40f90933
00112623
00912223
40295913
02090063
00000413
00000493
00042783
00148493
00440413
000780e7
fe9918e3
00000793
00000913
40f90933
40295913
02090063
00000413
00000493
00042783
00148493
00440413
000780e7
fe9918e3
00c12083
00812403
00412483
00012903
01010113
00008067
00f00313
00050713
02c37e63
00f77793
0a079063
08059263
ff067693
00f67613
00e686b3
00b72023
00b72223
00b72423
00b72623
01070713
fed766e3
00061463
00008067
40c306b3
00269693
00000297
005686b3
00c68067
00b70723
00b706a3
00b70623
00b705a3
00b70523
00b704a3
00b70423
00b703a3
00b70323
00b702a3
00b70223
00b701a3
00b70123
00b700a3
00b70023
00008067
0ff5f593
00859693
00d5e5b3
01059693
00d5e5b3
f6dff06f
00279693
00000297
005686b3
00008293
fa0680e7
00028093
ff078793
40f70733
00f60633
f6c378e3
f3dff06f
fd010113
01412c23
59402a03
03212023
02112623
148a2903
02812423
02912223
01312e23
01512a23
01612823
01712623
01812423
04090063
00050b13
00058b93
00100a93
fff00993
00492483
fff48413
02044263
00249493
009904b3
040b8463
1044a783
05778063
fff40413
ffc48493
ff3416e3
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
00492783
0044a683
fff78793
04878e63
0004a223
fa0688e3
18892783
008a9733
00492c03
00f777b3
02079263
000680e7
00492703
148a2783
01871463
f92784e3
f80788e3
00078913
f5dff06f
18c92783
0844a583
00f77733
00071c63
000b0513
000680e7
fcdff06f
00892223
fa9ff06f
00058513
000680e7
fb9ff06f
ff010113
00812423
00000793
00000413
40f40433
00912223
00112623
40245493
02048063
ffc40413
00f40433
00042783
fff48493
ffc40413
000780e7
fe0498e3
00c12083
00812403
00412483
01010113
00008067
00050593
00000693
00000613
00000513
0040006f
59402703
14872783
04078c63
0047a703
01f00813
06e84e63
00271813
02050663
01078333
08c32423
1887a883
00100613
00e61633
00c8e8b3
1917a423
10d32423
00200693
02d50463
00170713
00e7a223
010787b3
00b7a423
00000513
00008067
14c70793
14f72423
fa5ff06f
18c7a683
00170713
00e7a223
00c6e6b3
18d7a623
010787b3
00b7a423
00000513
00008067
fff00513
00008067
05d00893
00000073
00054463
0000006f
ff010113
00812423
00050413
00112623
40800433
00c000ef
00852023
0000006f
200007b7
4307a503
00008067
00000793
00078663
44400513
f0dff06f
00008067
20000000
00000000
200002ec
20000354
200003bc
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000001
00000000
abcd330e
e66d1234
0005deec
0000000b
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
20000000
00000054
0000009c
00000580
