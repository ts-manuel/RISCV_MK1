00026197
97018193
08000117
ff810113
00022297
65028293
04000317
fe830313
04001397
9d438393
406383b3
00038e63
0002ae03
01c32023
00428293
00430313
ffc38393
fe9ff06f
04001297
a6028293
04259317
b0430313
40530333
00030a63
0002a023
00428293
ffc30313
ff1ff06f
0040006f
00026197
8fc18193
04001517
97850513
04259617
ad060613
40a60633
00000593
64c020ef
00016517
6ec50513
00050863
00009517
cb050513
6d8160ef
5cd010ef
00012503
00410593
00000613
340220ef
0e40106f
ff010113
00812423
04001437
aa844783
00112623
02079263
00000793
00078a63
04001537
9f450513
00000097
000000e7
00100793
aaf40423
00c12083
00812403
01010113
00008067
00000793
00078e63
040015b7
04001537
aac58593
9f450513
00000317
00000067
00008067
04259737
b0c72783
00078a63
00a78533
b0a72623
00078513
00008067
042597b7
b5478793
00a78533
b0a72623
00078513
00008067
04259737
b2070ea3
04259737
00100793
b2070e23
04001737
9ef700a3
04001737
9ef70023
00008067
0f10206f
040017b7
9dc7a783
1207c063
04001837
00379713
9e184683
040017b7
fe010113
ac478793
00e787b3
00112e23
00812c23
00912a23
01212823
01312623
01412423
0007a703
10069a63
0047a783
04259937
b3892483
00f70733
0c976a63
200007b7
1047c983
0c098a63
042597b7
b2c7da03
042597b7
b347d403
003a5513
00040593
6bd000ef
00800793
00050593
18fa0263
00100793
1ef40463
00048713
00000693
ffff8637
200008b7
00374783
00174403
00274503
00074803
00879793
00841413
00a7e7b3
01046433
00c787b3
00c40433
01079793
01041413
0107d793
00f46433
1088a023
00168693
00b70733
fad99ee3
00098513
649000ef
00a484b3
b2992c23
200007b7
01c12083
1087a023
01812403
01412483
01012903
00c12983
00812a03
02010113
00008067
00008067
042597b7
b2092c23
b2078ea3
01c12083
01812403
01412483
01012903
00c12983
00812a03
02010113
00008067
01974503
01874e03
01a74783
01774583
01b74603
02374683
01674303
00851513
02274883
01c56533
01079793
00a7e7b3
00859593
01861613
0065e5b3
00f66633
00869693
042597b7
0116e6b3
b2b79a23
00025537
042597b7
04259437
02870713
b2d79623
d0850513
042597b7
b2c42823
b2e7ac23
9e0800a3
4a0020ef
b3042583
05f5e537
10050513
589000ef
01c12083
01812403
01051513
200007b7
10a7a223
01412483
01012903
00c12983
00812a03
02010113
00008067
00100793
02f40c63
00048793
00000693
20000637
0007c403
0017c703
00168693
01841413
00871713
00e46433
10862023
00b787b3
fed990e3
ea9ff06f
00048713
00000793
20000637
00074403
00178793
00b70733
00841693
01841413
00d46433
10862023
fef992e3
e79ff06f
00048793
00000713
ffff8537
20000637
0017c403
0007c683
00170713
00841413
00d46433
00a40433
01041693
0106d693
01041413
00d46433
10862023
00b787b3
fce998e3
e31ff06f
fb010113
04812423
00025437
d2c40593
04112623
04912223
05212023
03312e23
03412c23
03512a23
000103a3
00012623
435020ef
0a050263
00100a13
06400913
000259b7
07300493
00025ab7
0240006f
00050593
d34a8513
354020ef
00000a13
d2c40593
00000513
3fd020ef
02050863
00054783
05278863
fc979ce3
d3098593
00c10613
00250513
610020ef
d2c40593
00000513
3d1020ef
fc051ce3
020a1e63
04c12083
04812403
04412483
04012903
03c12983
03812a03
03412a83
05010113
00008067
00710613
d3098593
00250513
5c8020ef
f8dff06f
00c12583
fc0582e3
00714603
00025537
d5850513
2c0020ef
00714583
00400793
22b7e063
04001937
00359793
ac490913
00f907b3
0007a503
1b1010ef
00c12403
00714483
00040513
191010ef
00349793
00f907b3
00a7a023
0087a223
20050463
00000a93
08040463
00023a37
000239b7
06600493
108a0a13
2a498993
000a8513
175000ef
225000ef
14a4e463
00251793
014787b3
0007a783
00078067
00451513
0f057413
205000ef
02a4e063
00251793
013787b3
0007a783
00078067
008507b3
fd078793
0ff7f413
00714783
00379793
00f907b3
0007a783
015787b3
00878023
00c12783
001a8a93
f8faeae3
000257b7
ddc78793
0087a683
00c7a703
0007a583
0047a603
0107d783
02d12223
02e12423
02f11623
676f77b7
25078793
00f12823
737367b7
57278793
00f12a23
005b27b7
03a78793
00f12c23
000067b7
d2578793
00f11423
00b12e23
02c12023
00010523
01c10713
02000793
200006b7
00f68023
00174783
00170713
fe079ae3
01014783
01010713
200006b7
00078a63
00f68023
00174783
00170713
fe079ae3
200007b7
03100713
00e78023
03000713
00e78023
00e78023
00814783
00810713
200006b7
00078a63
00f68023
00174783
00170713
fe079ae3
00a00513
164020ef
dfdff06f
00000413
ed1ff06f
00f40413
0ff47413
ee9ff06f
00e40413
0ff47413
eddff06f
0f000413
eb1ff06f
0e000413
ea9ff06f
0d000413
ea1ff06f
0c000413
e99ff06f
00d40413
0ff47413
eb1ff06f
00c40413
0ff47413
ea5ff06f
00b40413
0ff47413
e99ff06f
00a40413
0ff47413
e8dff06f
00025537
00400613
d7c50513
088020ef
d79ff06f
0a000413
e4dff06f
0b000413
e45ff06f
00025537
00400613
00048593
da850513
060020ef
d51ff06f
06600793
02a7e463
00023737
00251793
44070713
00e787b3
0007a783
00078067
fd050513
0ff57513
00008067
00000513
00008067
00c00513
00008067
00f00513
00008067
00d00513
00008067
00e00513
00008067
00a00513
00008067
00b00513
00008067
000257b7
ddc78793
0087a683
00c7a703
0007a583
0047a603
0107d783
fb010113
04912223
02f11623
676f77b7
25078793
00f12823
737367b7
57278793
00f12a23
005b27b7
03a78793
00f12c23
000067b7
d2578793
02d12223
02e12423
00f11623
04112623
04812423
05212023
03312e23
00050493
00b12e23
02c12023
00010723
01c10713
02000793
200006b7
00f68023
00174783
00170713
fe079ae3
01014783
01010713
200006b7
00078a63
00f68023
00174783
00170713
fe079ae3
00a00593
00048513
0a5000ef
00900793
03050413
0497ce63
02000713
02000513
200007b7
00a78023
00e78023
0ff47413
00878023
00c14783
00c10713
200006b7
00078a63
00f68023
00174783
00170713
fe079ae3
04c12083
04812403
04412483
04012903
03c12983
05010113
00008067
00a00593
00048513
7b0000ef
00a00593
00050993
7a4000ef
00050913
00a00593
00098513
019000ef
03050713
06300793
0ff77713
0097d863
03090513
0ff57513
f71ff06f
02000513
f69ff06f
042597b7
b3d7c783
00078463
801ff06f
00008067
042597b7
b3c7c503
04050863
04001737
9d872703
04074263
04001637
00371693
9e064803
04001737
ac470713
00d70733
00072683
02081463
00472703
04259eb7
b20eae03
00e686b3
07c6fe63
b20ea023
b2078e23
00008067
00008067
040017b7
04259737
ae478793
b2f72423
0412d7b7
04259737
ae478793
b2f72223
042597b7
b2d7a023
00025537
042597b7
ff010113
b007ae23
df050513
042597b7
00112623
b007ac23
9e060023
03c020ef
00c12083
200007b7
32200713
20e7a423
01010113
00008067
04259637
b1462783
00013737
bff70713
16f74863
20000737
20472703
040016b7
9d46c883
01071593
0105d593
2e089a63
000106b7
ff068693
00d77733
042592b7
2c071c63
00700713
06b75263
042598b7
b288a703
200006b7
10078793
00072f03
02070313
ff858593
21e6a023
00472f03
21e6a023
00872f03
21e6a023
00c72f03
21e6a023
01072f03
21e6a023
01472f03
21e6a023
01872f03
21e6a023
01c72703
b268a423
20e6a023
b0f62a23
00300713
04b75063
042595b7
b285a703
200006b7
08078793
00072303
01070893
2066a023
00472303
2066a023
00872303
2066a023
00c72703
b315a423
20e6a023
b0f62a23
b102af83
000137b7
bff78793
e9f7cce3
042593b7
b243a683
00050893
00000793
0006a023
00100313
13f00f13
000e4603
001e0e13
02060e63
16089e63
00f605b3
01f7f713
0006a603
00e31733
00178793
00e66733
00e6a023
01f7f713
00071863
0006a223
00050813
00468693
fcf59ce3
0018c893
faff5ce3
b3cea023
00080463
b2d3a223
140f8f93
b1f2a823
00008067
042595b7
b185a703
042598b7
00200693
00170793
b0f5ac23
b1c8a783
12e6c663
04001737
ae470713
042592b7
00279693
00f686b3
00469793
40d787b3
00e79793
00f70733
042597b7
b2e7a423
040016b7
00100793
9cf68a23
200007b7
2047a703
b0062a23
000107b7
00f77733
f00702e3
200007b7
2007a223
b1462783
9c068a23
03000593
042598b7
b288a703
200006b7
20078793
00072f03
04070313
21e6a023
00472f03
21e6a023
00872f03
21e6a023
00c72f03
21e6a023
01072f03
21e6a023
01472f03
21e6a023
01872f03
21e6a023
01c72f03
21e6a023
02072f03
21e6a023
02472f03
21e6a023
02872f03
21e6a023
02c72f03
21e6a023
03072f03
21e6a023
03472f03
21e6a023
03872f03
21e6a023
b268a423
03c72703
20e6a023
b0f62a23
da5ff06f
00f60633
00178793
01f7f713
00071863
0006a223
00088813
00468693
fec794e3
e9dff06f
00279713
00f70733
00178793
01f7d313
00471693
40e686b3
006787b3
04001737
00e69693
ae470713
0017f793
406787b3
00d706b3
042592b7
04259337
b2d32223
b0f8ae23
b002a823
b005ac23
e99ff06f
ff058593
ee9ff06f
042592b7
ec1ff06f
fd010113
03212023
00025937
02912223
01512a23
fff00793
04001ab7
040014b7
d2c90593
02112623
02812423
01312e23
01412c23
01612823
01712623
9cfaae23
9cf4ac23
2f0020ef
0a050c63
00050793
00100b13
06100a13
00025437
07600993
00025bb7
0280006f
00078593
e1cb8513
20d010ef
00000b13
d2c90593
00000513
2b4020ef
00050793
02050a63
0007c703
05470e63
9d848613
d3040593
00278513
fd3714e3
4c5010ef
d2c90593
00000513
284020ef
00050793
fc051ae3
040b1263
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
03010113
00008067
9dca8613
d3040593
00278513
471010ef
f7dff06f
9d84a603
9dcaa583
00025537
e4050513
16d010ef
00100793
04259737
b2f70ea3
04259737
b2f70e23
04001737
9ef700a3
04001737
9ef70023
ad4ff0ef
02812403
02c12083
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
03010113
ab1ff06f
00500793
02a7e663
000237b7
00f5f593
5dc78793
00b787b3
0007c703
020007b7
00278793
00f50533
00451513
00e52023
00008067
000237b7
5dc78793
00f57693
00455713
00d786b3
00855593
00f77713
00e78733
0006c883
00c55613
00f5f593
00074803
00b785b3
01055693
00f67613
20000737
00c78633
0005c583
00f6f693
01455513
03172023
00d786b3
00064603
00f57513
03072823
0006c683
00a787b3
04b72023
0007c783
04c72823
06d72023
06f72823
00008067
042597b7
b3e7c703
00100513
02071063
20000737
00072703
042596b7
00f75513
00157513
b2e68fa3
b2a78f23
00008067
04259737
b3e74783
00078a63
042597b7
b3f7c503
b2070f23
00008067
042595b7
20000637
000086b7
00062783
0ff7f513
b2a58fa3
00d7f7b3
fe0788e3
fd9ff06f
20000737
00472783
0107d793
fe078ce3
00a70023
00008067
00060513
02c05463
00c58833
20000737
0005c683
00158593
00472783
0107d793
fe078ce3
00d70023
feb814e3
00008067
00060513
06c05463
04259637
b3e64783
00a58333
042596b7
200008b7
00008837
0140006f
b3f6c703
fee58fa3
00000793
02658c63
00158593
fe0796e3
0008a783
0ff7f713
b2e68fa3
0107f7b3
fc079ee3
0008a783
0ff7f713
b2e68fa3
0107f7b3
fc078ee3
fc5ff06f
b2060f23
00008067
00050613
00000513
0015f693
00068463
00c50533
0015d593
00161613
fe0596e3
00008067
06054063
0605c663
00058613
00050593
fff00513
02060c63
00100693
00b67a63
00c05863
00161613
00169693
feb66ae3
00000513
00c5e663
40c585b3
00d56533
0016d693
00165613
fe0696e3
00008067
00008293
fb5ff0ef
00058513
00028067
40a00533
00b04863
40b005b3
f9dff06f
40b005b3
00008293
f91ff0ef
40a00533
00028067
00008293
0005ca63
00054c63
f79ff0ef
00058513
00028067
40b005b3
fe0558e3
40a00533
f61ff0ef
40b00533
00028067
ff010113
00000593
00812423
00112623
00050413
0f5070ef
000257b7
0d07a503
03c52783
00078463
000780e7
00040513
0111a0ef
00c59783
fe010113
00812c23
01312623
00112e23
00912a23
01212823
0087f693
00058413
00050993
10069c63
00001737
80070713
0045a683
00e7e7b3
00f59623
18d05663
02842703
0c070c63
01079793
0107d793
000016b7
0009a483
00d7f6b3
0009a023
01c42583
16069863
00100693
00000613
00098513
000700e7
fff00793
18f50e63
00c45783
02842703
01c42583
0047f793
00078e63
00442683
03042783
40d50533
00078663
03c42783
40f50533
00050613
00000693
00098513
000700e7
fff00793
10f51e63
0009a703
00c41783
16070a63
01d00693
00d70663
01600693
0cd71463
01042683
fffff737
7ff70713
00e7f7b3
00f41623
00042223
00d42023
03042583
0099a023
00058c63
04040793
00f58663
00098513
71c000ef
02042823
00000513
01c12083
01812403
01412483
01012903
00c12983
02010113
00008067
0105a903
fc090ee3
0005a483
01079713
01075713
00377713
0125a023
412484b3
00000793
00071463
0145a783
00f42423
00904863
fadff06f
00a90933
fa9052e3
02442783
01c42583
00048693
00090613
00098513
000780e7
40a484b3
fca04ee3
00c45783
fff00513
0407e793
01c12083
00f41623
01812403
01412483
01012903
00c12983
02010113
00008067
03c5a703
e6e04ae3
f4dff06f
05042503
eb5ff06f
00c45783
fffff737
7ff70713
00e7f7b3
01042683
01079793
4107d793
00c7d713
00f41623
00042223
00d42023
00177793
ee0788e3
04a42823
ee9ff06f
0009a783
e60782e3
01d00713
02e78863
01600713
02e78463
00c45783
0407e793
00f41623
ee5ff06f
fffff737
7ff70713
01042683
00e7f7b3
fa9ff06f
0099a023
00000513
ec5ff06f
fe010113
00812c23
00112e23
00050413
00050663
03852783
02078063
00c59783
02079663
01c12083
01812403
00000513
02010113
00008067
00b12623
40c000ef
00c12583
00c59783
fc078ee3
00040513
01812403
01c12083
02010113
d41ff06f
06050863
fe010113
040017b7
00812c23
00050413
9e47a503
00112e23
00050663
03852783
02078a63
00c41783
00079c63
01c12083
01812403
00000513
02010113
00008067
00040593
01812403
01c12083
02010113
ce9ff06f
00a12623
38c000ef
00c41783
00c12503
fc0784e3
fd9ff06f
000257b7
0d07a503
000015b7
44058593
0a90006f
00000513
00008067
000095b7
c3458593
0950006f
00000513
00008067
fe010113
000017b7
00112e23
00812c23
00912a23
01212823
01312623
01412423
01512223
01612023
00452403
52c78793
02f52e23
2ec50713
00300793
2ee52423
2ef52223
2e052023
00400793
00050913
00f42623
00800613
00000593
06042223
00042023
00042223
00042423
00042823
00042a23
00042c23
05c40513
124010ef
00003b37
00892483
00003ab7
00003a37
000039b7
c18b0b13
c7ca8a93
d04a0a13
d6c98993
000107b7
03642023
03542223
03442423
03342623
00842e23
00978793
00f4a623
00800613
00000593
0604a223
0004a023
0004a223
0004a423
0004a823
0004aa23
0004ac23
05c48513
0b4010ef
00c92403
000207b7
0364a023
0354a223
0344a423
0334a623
0094ae23
01278793
00f42623
06042223
00042023
00042223
00042423
00042823
00042a23
00042c23
05c40513
00800613
00000593
064010ef
01c12083
03642023
03542223
03442423
03342623
00842e23
01812403
00100793
02f92c23
01412483
01012903
00c12983
00812a03
00412a83
00012b03
02010113
00008067
ff010113
fff58793
00812423
00179413
00f40433
00241413
00f40433
00341413
01212023
00058913
07440593
00912223
00112623
031000ef
00050493
02050063
00c50513
0004a023
0124a223
00a4a423
06840613
00000593
7c5000ef
00c12083
00812403
00012903
00048513
00412483
01010113
00008067
fe010113
000257b7
01212823
0d07a903
01312623
00112e23
03892783
00812c23
00912a23
01412423
00050993
0a078a63
2e090913
fff00493
00400a13
00492783
00892403
fff78793
0007d863
0840006f
06840413
06978e63
00c41703
fff78793
fe0718e3
ffff07b7
00178793
06042223
00042023
00042223
00042423
00f42623
00042823
00042a23
00042c23
00800613
00000593
05c40513
70d000ef
02042823
02042a23
04042223
04042423
01c12083
00040513
01812403
01412483
01012903
00c12983
00812a03
02010113
00008067
00092403
00040c63
00040913
f61ff06f
00090513
d21ff0ef
f49ff06f
1ac00593
00098513
6f8000ef
00050413
02050663
00c50513
00042023
01442223
00a42423
1a000613
00000593
68d000ef
00892023
00040913
f19ff06f
00092023
00c00793
00f9a023
f79ff06f
000257b7
0d07a503
000095b7
c3458593
5440006f
03852783
00078463
00008067
cadff06f
00008067
00008067
00008067
00008067
040017b7
9e47a503
000015b7
52458593
46c0006f
040017b7
9e47a503
000015b7
53858593
4580006f
fe010113
01312623
040009b7
00812c23
00912a23
01212823
01412423
00112e23
00058a13
00050913
44898993
6c1000ef
0089a703
000017b7
fef78413
00472483
41440433
ffc4f493
00940433
00c45413
fff40413
00c41413
00f44e63
00000593
00090513
15c010ef
0089a783
009787b3
02f50863
00090513
679000ef
01c12083
01812403
01412483
01012903
00c12983
00812a03
00000513
02010113
00008067
408005b3
00090513
118010ef
fff00793
04f50a63
042597b7
ae478793
0007a703
0089a683
408484b3
0014e493
40870733
00090513
0096a223
00e7a023
615000ef
01c12083
01812403
01412483
01012903
00c12983
00812a03
00100513
02010113
00008067
00000593
00090513
0b4010ef
0089a703
00f00693
40e507b3
f4f6dce3
040016b7
9e86a683
0017e793
00f72223
40d50533
042596b7
aea6a223
f39ff06f
12058a63
ff010113
00812423
00912223
00058413
00050493
00112623
591000ef
ffc42803
ff840713
040005b7
ffe87793
00f70633
44858593
00462683
0085a503
ffc6f693
1ac50a63
00d62223
00187813
00d60533
0a081063
ff842303
00452803
04000537
40670733
00872883
45050513
006787b3
00187813
14a88063
00c72303
0068a623
01132423
1e080463
0017e693
00d72223
00f62023
1ff00693
0af6e863
ff87f693
00868693
0045a503
00d586b3
0006a603
0057d813
00100793
010797b3
00a7e7b3
ff868513
00a72623
00c72423
00f5a223
00e6a023
00e62623
00812403
00c12083
00048513
00412483
01010113
4c10006f
00452503
00157513
02051e63
04000537
00d787b3
45050513
00862683
0017e893
00f70833
16a68863
00c62603
00c6a623
00d62423
01172223
00f82023
f69ff06f
00008067
0017e693
fed42e23
00f62023
1ff00693
f4f6fce3
0097d693
00400613
0ed66c63
0067d693
03968813
03868613
00381813
01058833
00082683
ff880813
12d80863
0046a603
ffc67613
00c7f663
0086a683
fed818e3
00c6a803
01072623
00d72423
00812403
00c12083
00e82423
00048513
00412483
00e6a623
01010113
3fd0006f
14081663
00c62583
00862603
00f686b3
00812403
00b62623
00c5a423
0016e793
00c12083
00f72223
00048513
00d70733
00412483
00d72023
01010113
3bd0006f
00187813
00d786b3
02081063
ff842503
40a70733
00c72783
00872603
00a686b3
00f62623
00c7a423
040017b7
0016e613
9ec7a783
00c72223
00e5a423
eaf6e4e3
042597b7
b487a583
00048513
c7dff0ef
e95ff06f
01400613
02d67463
05400613
06d66463
00c7d693
06f68813
06e68613
00381813
efdff06f
00d787b3
e99ff06f
05c68813
05b68613
00381813
ee5ff06f
00e5aa23
00e5a823
00a72623
00a72423
01172223
00f82023
e3dff06f
0045a503
40265613
00100793
00c797b3
00a7e7b3
00f5a223
ed5ff06f
15400613
00d66c63
00f7d693
07868813
07768613
00381813
e91ff06f
55400613
00d66c63
0127d693
07d68813
07c68613
00381813
e75ff06f
3f800813
07e00613
e69ff06f
0017e693
00d72223
00f62023
dcdff06f
fe010113
01212823
01312623
01412423
01512223
01612023
00112e23
00812c23
00912a23
00058b13
2e050a93
00000a13
00100993
fff00913
004aa483
008aa403
fff48493
0204c663
00c45783
fff48493
00f9fc63
00e41783
00040513
01278663
000b00e7
00aa6a33
06840413
fd249ee3
000aaa83
fc0a92e3
01c12083
01812403
01412483
01012903
00c12983
00412a83
00012b03
000a0513
00812a03
02010113
00008067
fd010113
03212023
01312e23
01412c23
01512a23
01612823
01712623
02112623
02812423
02912223
00050a93
00058b93
2e050b13
00000a13
00100993
fff00913
004b2483
008b2403
fff48493
0204c863
00c45783
fff48493
00f9fe63
00e41783
00040593
000a8513
01278663
000b80e7
00aa6a33
06840413
fd249ce3
000b2b03
fc0b10e3
02c12083
02812403
02412483
02012903
01c12983
01412a83
01012b03
00c12b83
000a0513
01812a03
03010113
00008067
ff010113
00812423
01212023
00000793
00000913
40f90933
00112623
00912223
40295913
02090063
00000413
00000493
00042783
00148493
00440413
000780e7
fe9918e3
00000793
00000913
40f90933
40295913
02090063
00000413
00000493
00042783
00148493
00440413
000780e7
fe9918e3
00c12083
00812403
00412483
00012903
01010113
00008067
040017b7
00050593
9e47a503
0140006f
040017b7
00050593
9e47a503
aedff06f
fd010113
01312e23
02112623
02812423
02912223
03212023
01412c23
01512a23
01612823
01712623
01812423
01912223
00b58793
01600713
00050993
06f76663
01000793
1eb7e663
04d000ef
01000493
01800793
00200613
04000937
44890913
00f907b3
0047a403
ff878713
20e40a63
00442783
00c42683
00842603
ffc7f793
00f407b3
0047a703
00d62623
00c6a423
00176713
00098513
00e7a223
7fc000ef
00840513
1980006f
ff87f493
1807c263
18b4e063
7e0000ef
1f700793
4697f663
0094d793
1a078663
00400713
3cf76c63
0064d793
03978613
03878513
00361693
04000937
44890913
00d906b3
0046a403
ff868693
02868663
00f00593
0100006f
32075c63
00c42403
00868c63
00442783
ffc7f793
40978733
fee5d4e3
00050613
01092403
00890893
17140863
00442583
00f00713
ffc5f593
409587b3
40f74c63
01192a23
01192823
3e07d663
1ff00793
2eb7ea63
ff85f793
00878793
00492503
00f907b3
0007a683
0055d593
00100713
00b71733
00a76733
ff878593
00b42623
00d42423
00e92223
0087a023
0086a623
40265793
00100593
00f595b3
10b76863
00e5f7b3
02079463
00159593
ffc67613
00e5f7b3
00460613
00079a63
00159593
00e5f7b3
00460613
fe078ae3
00f00813
00361313
00690333
00030513
00c52783
00060e13
2ef50263
0047a703
00078413
00c7a783
ffc77713
409706b3
2ed84263
fe06c2e3
00e40733
00472683
00842603
00098513
0016e693
00d72223
00f62623
00c7a423
674000ef
00840513
0100006f
00c00793
00f9a023
00000513
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
03010113
00008067
20000693
04000613
03f00513
e65ff06f
00c7a403
00260613
de8794e3
01092403
00890893
e9141ce3
00492703
40265793
00100593
00f595b3
eeb77ce3
00892403
00442b03
ffcb7b13
009b6863
409b07b3
00f00713
14f74663
042597b7
04001cb7
b487aa83
9e8ca703
fff00793
01640a33
01548ab3
34f70a63
000017b7
00f78793
00fa8ab3
fffff7b7
00fafab3
000a8593
00098513
065000ef
fff00793
00050b93
28f50c63
29456863
04259c37
ae4c0c13
000c2583
00ba85b3
00bc2023
00058793
3aaa0463
9e8ca683
fff00713
3ae68c63
414b8a33
00fa07b3
00fc2023
007bfc93
300c8663
000017b7
419b8bb3
00878593
008b8b93
419585b3
015b8ab3
fff78793
415585b3
00f5fa33
000a0593
00098513
7e8000ef
fff00793
3cf50063
41750533
01450ab3
000c2783
01792423
001aea93
00fa05b3
00bc2023
015ba223
35240863
00f00693
3566f863
00442703
ff4b0793
ff87f793
00177713
00f76733
00e42223
00500613
00f40733
00c72223
00c72423
36f6ee63
004baa83
000b8413
042597b7
b447a703
00b77463
b4b7a223
042597b7
b407a703
1ab77663
b4b7a023
1a40006f
0014e713
00e42223
009404b3
00992423
0017e793
00098513
00f4a223
46c000ef
00840513
e09ff06f
00c42683
00842603
c41ff06f
0095d793
00400713
14f77263
01400713
22f76a63
05c78693
05b78713
00369693
00d906b3
0006a783
ff868693
1cf68863
0047a703
ffc77713
00e5f663
0087a783
fef698e3
00c7a683
00492703
00d42623
00f42423
0086a423
0087a623
cf1ff06f
01400713
12f77663
05400713
1ef76a63
00c4d793
06f78613
06e78513
00361693
c1dff06f
001e0e13
003e7793
00850513
10078e63
00c52783
d09ff06f
00842603
0014e593
00b42223
00f62623
00c7a423
009404b3
00992a23
00992823
0016e793
0114a623
0114a423
00f4a223
00e40733
00098513
00d72023
37c000ef
00840513
d19ff06f
0034d613
00848793
b29ff06f
00b405b3
0045a783
00098513
0017e793
00f5a223
350000ef
00840513
cedff06f
0014e713
00e42223
009404b3
00992a23
00992823
0017e713
0114a623
0114a423
00e4a223
00b405b3
00098513
00f5a023
314000ef
00840513
cb1ff06f
0065d793
03978693
03878713
00369693
ec5ff06f
11240e63
00892403
00442a83
ffcafa93
409a87b3
009ae663
00f00713
e4f748e3
00098513
2d0000ef
00000513
c6dff06f
05c78613
05b78513
00361693
b01ff06f
00832783
fff60613
1c679263
00367793
ff830313
fe0796e3
00492703
fff5c793
00e7f7b3
00f92223
00159593
c8b7eee3
c8058ce3
00f5f733
00071a63
00159593
00f5f733
004e0e13
fe070ae3
000e0613
b9dff06f
010a8a93
cc1ff06f
00492503
40275593
00100713
00b71733
00a76733
00e92223
e39ff06f
015b85b3
40b005b3
01459593
0145da13
000a0593
00098513
4f4000ef
fff00793
d0f518e3
00000a13
d11ff06f
05400713
08f76263
00c5d793
06f78693
06e78713
00369693
dc5ff06f
15400713
08f76263
00f4d793
07878613
07778513
00361693
a25ff06f
04259c37
ae4c0c13
000c2783
00fa87b3
00fc2023
c61ff06f
014a1713
c4071ce3
00892403
015b0ab3
001aea93
01542223
cfdff06f
9f7ca423
c55ff06f
000b8413
cedff06f
00100793
00fba223
eb9ff06f
15400713
06f76263
00f5d793
07878693
07778713
00369693
d3dff06f
55400713
06f76263
0124d793
07d78613
07c78513
00361693
99dff06f
ff8c8c93
019a8ab3
417a8ab3
00000a13
c3dff06f
00840593
00098513
b84ff0ef
00892403
000c2583
00442a83
c79ff06f
55400713
02f76463
0125d793
07d78693
07c78713
00369693
cd5ff06f
3f800693
07f00613
07e00513
941ff06f
3f800693
07e00713
cb9ff06f
00492783
e59ff06f
00f00313
00050713
02c37e63
00f77793
0a079063
08059263
ff067693
00f67613
00e686b3
00b72023
00b72223
00b72423
00b72623
01070713
fed766e3
00061463
00008067
40c306b3
00269693
00000297
005686b3
00c68067
00b70723
00b706a3
00b70623
00b705a3
00b70523
00b704a3
00b70423
00b703a3
00b70323
00b702a3
00b70223
00b701a3
00b70123
00b700a3
00b70023
00008067
0ff5f593
00859693
00d5e5b3
01059693
00d5e5b3
f6dff06f
00279693
00000297
005686b3
00008293
fa0680e7
00028093
ff078793
40f70733
00f60633
f6c378e3
f3dff06f
00008067
00008067
fc010113
02c12423
02d12623
02e12823
02f12a23
03012c23
03112e23
00058613
00852583
02810693
00112e23
00d12623
618030ef
01c12083
04010113
00008067
04001337
9e432303
fc010113
02c12423
02d12623
02b12223
02e12823
02f12a23
03012c23
03112e23
00832583
02410693
00050613
00030513
00112e23
00d12623
5c8030ef
01c12083
04010113
00008067
00852603
01c0006f
040017b7
9e47a783
00050593
0087a603
00078513
0040006f
fe010113
01212c23
00112e23
00050913
00050663
03852783
04078663
00862783
fff78793
00f62423
0007dc63
01862703
04e7c663
0ff5f793
00a00713
04e78063
00062783
0ff5f513
00178713
00e62023
00b78023
01c12083
01812903
02010113
00008067
00c12623
00b12423
fa9fe0ef
00c12603
00812583
fa5ff06f
01c12083
00090513
01812903
02010113
6390506f
ff010113
040017b7
01212023
9e47a903
00812423
00912223
00112623
00050493
00058413
00090663
03892783
04078a63
00842783
fff78793
00f42423
0007dc63
01842703
04e7c463
0ff4f793
00a00713
02e78e63
00042783
0ff4f513
00178713
00e42023
00978023
00c12083
00812403
00412483
00012903
01010113
00008067
00090513
f01fe0ef
fa9ff06f
00040613
00812403
00c12083
00048593
00090513
00412483
00012903
01010113
5890506f
fc010113
02812c23
00050413
00058513
02912a23
02112e23
00058493
660000ef
000257b7
e6878793
02f12423
00100793
02f12623
03842703
02010793
00150693
00f12a23
00200793
02912023
02a12223
00d12e23
00f12c23
00842583
04070e63
00c59783
01279713
02074263
0645a703
000026b7
00d7e7b3
ffffe6b7
fff68693
00d77733
00f59623
06e5a223
01410613
00040513
360060ef
03c12083
03812403
00a03533
40a00533
03412483
00a56513
04010113
00008067
00040513
00b12623
e15fe0ef
00c12583
f99ff06f
040017b7
00050593
9e47a503
f29ff06f
ff010113
00812423
00912223
00050413
042594b7
00058513
00112623
b404a823
e84fd0ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
f6010113
08f12a23
20400793
06112e23
06812c23
08c12423
00058413
08d12623
08e12823
09012c23
09112e23
00f11a23
00a12423
00a12c23
508000ef
00050793
04001737
00f12623
00f12e23
9e472503
000037b7
c7478793
08810693
02f12423
00040613
00810593
fff00793
02012c23
04012623
00f11b23
00d12223
604000ef
07c12083
07812403
0a010113
00008067
f6010113
06812c23
08f12a23
00050413
20400793
00058513
06112e23
06912a23
08d12623
00060493
08e12823
09012c23
09112e23
00f11a23
00b12423
00b12c23
470000ef
00050793
00f12623
00f12e23
000037b7
c7478793
08c10693
02f12423
00048613
00810593
00040513
fff00793
02012c23
04012623
00f11b23
00d12223
570000ef
07c12083
07812403
07412483
0a010113
00008067
ff010113
00812423
00058413
00e59583
00112623
5090a0ef
02054063
05042783
00c12083
00a787b3
04f42823
00812403
01010113
00008067
00c45783
fffff737
fff70713
00e7f7b3
00c12083
00f41623
00812403
01010113
00008067
00000513
00008067
00c59783
fe010113
00812c23
00912a23
01212823
01312623
00112e23
1007f713
00058413
00050493
00060913
00068993
04071063
fffff737
fff70713
00e7f7b3
00e41583
00f41623
01812403
01c12083
00098693
00090613
00c12983
01012903
00048513
01412483
02010113
3f10506f
00e59583
00200693
00000613
21c090ef
00c41783
fb1ff06f
ff010113
00812423
00058413
00e59583
00112623
1fc090ef
fff00793
02f50463
00c45783
00001737
00c12083
00e7e7b3
04a42823
00f41623
00812403
01010113
00008067
00c45783
fffff737
fff70713
00e7f7b3
00c12083
00f41623
00812403
01010113
00008067
00e59583
6650506f
0ff5f693
00357793
0c068063
00078e63
00054783
0a078663
0ad78663
00150513
00357793
fe0796e3
0ff5f593
00859793
00f5e5b3
00052703
01059313
00b36333
feff0837
00e34633
eff80813
010607b3
010705b3
fff64613
fff74713
00c7f7b3
00e5f733
808088b7
00e7e7b3
08088893
0117f7b3
02079a63
00452703
00450513
00674633
010707b3
010605b3
fff74713
fff64613
00e7f7b3
00c5f733
00e7e7b3
0117f7b3
fc078ae3
00054783
00078a63
08f68663
00154783
00150513
fe079ae3
00000513
00008067
00078c63
00054783
fe078ae3
00150513
00357793
fe0798e3
00052703
feff0637
eff60613
00c707b3
808086b7
fff74713
00e7f7b3
08068693
00d7f7b3
02079063
00452703
00450513
00c707b3
fff74713
00e7f7b3
00d7f7b3
fe0784e3
00054783
f8078ee3
00154783
00150513
fe079ce3
00008067
00008067
00b56733
fff00393
00377713
10071063
7f7f87b7
f7f78793
00052603
0005a683
00f672b3
00f66333
00f282b3
0062e2b3
10729263
08d61663
00452603
0045a683
00f672b3
00f66333
00f282b3
0062e2b3
0c729e63
06d61663
00852603
0085a683
00f672b3
00f66333
00f282b3
0062e2b3
0c729863
04d61663
00c52603
00c5a683
00f672b3
00f66333
00f282b3
0062e2b3
0c729263
02d61663
01052603
0105a683
00f672b3
00f66333
00f282b3
0062e2b3
0a729c63
01450513
01458593
f4d60ee3
01061713
01069793
00f71e63
01065713
0106d793
40f70533
0ff57593
02059063
00008067
01075713
0107d793
40f70533
0ff57593
00059463
00008067
0ff77713
0ff7f793
40f70533
00008067
00054603
0005c683
00150513
00158593
00d61463
fe0616e3
40d60533
00008067
00450513
00458593
fcd61ce3
00000513
00008067
00850513
00858593
fcd612e3
00000513
00008067
00c50513
00c58593
fad618e3
00000513
00008067
01050513
01058593
f8d61ee3
00000513
00008067
00357793
00050713
04079c63
7f7f86b7
f7f68693
fff00593
00072603
00470713
00d677b3
00d787b3
00c7e7b3
00d7e7b3
feb784e3
ffc74683
40a707b3
04068463
ffd74683
02068c63
ffe74503
00a03533
00f50533
ffe50513
00008067
fa0688e3
00074783
00170713
00377693
fe0798e3
40a70733
fff70513
00008067
ffd78513
00008067
ffc78513
00008067
040017b7
9e47a603
00100693
05c60613
0040006f
06050863
00054803
00150893
00058793
0080006f
04e80263
0007c703
00178793
fe071ae3
04080e63
0008c683
00058793
00188893
0080006f
fe0708e3
0007c703
00178793
fee69ae3
00068e63
fe088fa3
01162023
00008067
02068a63
00088513
fa5ff06f
00000893
01162023
00008067
00062503
f80518e3
00000513
00008067
00062023
00000513
00008067
01162023
00050023
00008067
00100693
f65ff06f
ae010113
50812c23
4f812c23
4f912a23
50112e23
50912a23
51212823
51312623
51412423
51512223
51612023
4f712e23
4fa12823
4fb12623
52010413
00c59703
fffff7b7
b1078793
008787b3
fffff2b7
00d7a023
01271693
00510133
00058c93
00050c13
0206c263
0645a683
000025b7
00b76733
ffffe5b7
fff58593
00b6f6b3
00ec9623
06dca223
fffff6b7
00064703
fc068793
008786b3
b6e6ae23
00160b13
fffff7b7
00071463
7240206f
b8078693
b0478793
008787b3
0007a023
fffff7b7
b1c78793
008787b3
0007a023
fffff7b7
b0c78793
008787b3
0007a023
fffff7b7
00024637
b1878793
008787b3
c0160d13
00023637
0007a023
5ec60793
fffff637
b1460613
00860633
00f62023
fc068793
fffff6b7
b0068693
008787b3
008686b3
00000b93
00f6a023
000c8793
00000d93
000b8c93
00078b93
00ed06b3
0006c683
0086f693
10069263
02500693
04d71863
000b4683
00000a13
00000493
05500613
06800313
06c00513
fdb68793
0ff7f793
001b0593
22f66063
fffff737
b1470713
00870733
00072703
00279793
00e787b3
0007a783
00078067
00058b13
004ba703
14e05663
000ba703
fffb4683
00074603
10d60263
fffff7b7
b1c78793
008787b3
0007a783
02078263
fffff7b7
b1c78793
008787b3
0007a783
0007aa03
000a0663
000a0513
bc5fe0ef
fffff7b7
b1878793
fffff2b7
008787b3
ae028293
0007a503
00540133
000012b7
00510133
51c12083
51812403
51412483
51012903
50c12983
50812a03
50412a83
50012b03
4fc12b83
4f812c03
4f412c83
4f012d03
4ec12d83
52010113
00008067
004ba703
02e05c63
000ba783
0007c703
00ed0733
00074703
00877713
02070863
004ba703
00178793
00fba023
fff70713
00eba223
001c8c93
fce048e3
000b8593
000c0513
0510d0ef
fc0500e3
000b4703
fffff7b7
fc078793
008786b3
b6e6ae23
001b0b13
e80716e3
f05ff06f
004ba683
00170713
00eba023
fff68713
00eba223
000b4703
fffff7b7
fc078793
008786b3
b6e6ae23
001c8c93
001b0b13
e4071ae3
ecdff06f
000b8593
000c0513
7e80d0ef
ea0506e3
000b8c93
fffff7b7
b1878793
008787b3
0007a783
00078863
00ccd783
0407f793
e8078ce3
fffff7b7
b1c78793
008787b3
0007a783
00079463
08d0206f
fffff7b7
b1c78793
008787b3
0007a783
0067d983
0007aa03
02098663
000a0493
00000913
0004a783
00448493
00190913
0007a503
a3dfe0ef
ffc4a783
0007a023
ff3912e3
fffff737
b1870713
fff00793
00870733
00f72023
e4dff06f
fffff7b7
b1c78793
008787b3
0007a783
e40782e3
0007aa03
e31ff06f
08fa7793
e00790e3
00249793
009784b3
00149493
00d484b3
fd048493
001b4683
00058b13
d95ff06f
00058b13
00400913
004ba703
3ce05063
040a7713
3c070863
00300713
64e902e3
00400713
1ae904e3
00100713
5ce90663
00200713
00e90463
0d00106f
00049463
fff00493
001a7993
010a7913
00099463
7740106f
00090463
0ec0206f
fffff7b7
b1078793
008787b3
0007a783
080a7313
00478993
0007aa03
00031463
2d80206f
f20a0ee3
08000513
939fe0ef
00050a93
ea050ce3
fffff7b7
b1c78793
008787b3
0007a683
00aa2023
0066d783
0046d703
00e7e463
3590106f
0006a503
00279713
00e50533
fffff737
b1c70713
00870733
00072703
00178793
01452023
00f71323
fffff7b7
b1078793
008787b3
0137a023
fffff7b7
afc78793
fffff737
008787b3
b0870713
0157a023
00870733
02000793
00f72023
000ba703
00074703
00ed0733
00074703
00877713
1c071c63
fffff737
fffff6b7
c9070313
b8870793
af468693
fc070713
00870733
008686b3
00e6a023
fc030713
00870333
fffff737
af870713
00870733
01472023
fffff737
fc078793
af070713
008787b3
00870733
01672023
00000993
000b8b13
00030a13
00090b93
00048913
00078493
7ac080ef
01351463
6650106f
fffff7b7
000b2703
af478793
008787b3
004b2683
0007a783
00074583
fff68693
01378633
00170713
00eb2023
c8b60823
00db2223
00300713
00198993
00ed9863
b887a783
00400713
00e78a63
00800613
00000593
00048513
f9dfe0ef
00098693
00048713
000a0613
000a8593
000c0513
291080ef
fff00693
00050d93
00d51463
5e10106f
00050463
0240206f
fffff7b7
aec78793
008787b3
000aa023
0137a023
2d9050ef
00050463
3b80206f
013c8cb3
fff90913
000b8463
30c0206f
fffff7b7
af878793
008787b3
0007a783
004a8a93
00079463
2f00206f
fffff7b7
afc78793
008787b3
0007a783
00000993
40fa8733
fffff7b7
b0878793
008787b3
0007a783
40275693
00f6e463
49c0206f
004b2703
00e04463
2d40206f
000b2703
00074703
00ed0733
00074703
00877713
00071463
ec0912e3
fffff7b7
af878793
008787b3
0007aa03
fffff7b7
af078793
008787b3
000b8913
000b0b93
0007ab03
ba091ee3
000aa023
020a0c63
fffff7b7
afc78793
008787b3
0007a783
40fa85b3
fffff7b7
b0878793
008787b3
0007a783
4025d713
00170713
00f77463
2340206f
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
b59ff06f
00fa7793
a60798e3
001b4683
002a6a13
00058b13
a15ff06f
00fa7793
c60788e3
a55ff06f
200a6a13
00011737
b0870793
fffff737
b0470713
00870733
00f72023
00058b13
01000793
fffff737
b0c70713
00870733
00f72023
004ba703
00300913
c4e044e3
000b8593
000c0513
3300d0ef
b40516e3
040a7713
c2071ce3
000ba683
0006c703
00ed0733
00074703
00877713
02071263
c1dff06f
00168693
00dba023
0006c783
00fd07b3
0007c783
0087f793
c00780e3
004ba783
001c8c93
fff78793
00fba223
fcf04ae3
000b8593
000c0513
2cc0d0ef
ae0514e3
000ba683
fc5ff06f
001a6a13
040a6a13
00058b13
00000913
bb1ff06f
001a6a13
00058b13
00200913
ba1ff06f
001a6a13
00011737
b0870793
fffff737
b0470713
00870733
00f72023
00058b13
00800793
f21ff06f
001a6a13
00010737
00058b13
36c70793
fffff737
b0470713
00870733
00f72023
00a00793
ef9ff06f
00fa7793
90079ee3
001b4683
00669463
5550106f
004a6a13
00058b13
8b9ff06f
00011737
00058b13
b0870793
fbdff06f
fffff7b7
b5078793
00878533
6880a0ef
00050b13
040a6a13
00100913
b01ff06f
00010737
36c70793
fffff737
b0470713
00870733
00f72023
fffff7b7
b0c78793
008787b3
00058b13
0007a023
00300913
acdff06f
00fa7793
88079ce3
001b4683
00a69463
4e10106f
001a6a13
00058b13
835ff06f
08fa7793
86079ce3
fffff7b7
b1c78793
008787b3
0007a783
00079463
5450106f
001b4683
080a6a13
00058b13
805ff06f
010a7713
00058b13
920712e3
fffff7b7
b1078793
008787b3
0007a783
008a7713
0007a683
00478613
00071463
6190106f
fffff7b7
b1078793
008787b3
01968023
00c7a023
8e9ff06f
220a6a13
db5ff06f
0144e4b3
fe049c63
001b4683
01000a13
00058b13
f9cff06f
00049463
fff00493
fffff6b7
afc68693
010a7793
008686b3
001a7713
00f6a023
00071463
7f90006f
00078463
2190106f
fffff7b7
b1078793
008787b3
0007a783
fffff6b7
af868693
0007a703
008686b3
00478793
00e6a023
fffff6b7
aec68693
008686b3
080a7313
00f6a023
00031463
5290106f
940708e3
08000513
b4cfe0ef
00050993
8c0506e3
fffff7b7
b1c78793
008787b3
fffff6b7
0007a783
af868693
008686b3
0006a683
0067d903
0047d703
00a6a023
00e96463
7940106f
0007a503
fffff7b7
b1c78793
008787b3
0007a783
00291713
00190913
01279323
fffff7b7
af878793
008787b3
0007a783
00e50533
fffff737
00f52023
fffff7b7
af078793
008787b3
af470713
0137a023
00870733
02000793
00f72023
fffff7b7
b8878a93
c5078793
00878a33
fc0a8793
00878ab3
fffff7b7
ae878793
008787b3
0167a023
fffff7b7
b0078793
008787b3
000a8b13
000a0a93
00048a13
0007a483
00000913
1ec080ef
fd250463
000ba703
004ba683
fffff537
00074583
fc050793
008787b3
01278633
00170713
fff68693
00eba023
c8b60823
00dba223
00300713
00190913
00ed9c63
b4050793
008787b3
0007a683
00400713
00e68a63
00800613
00000593
00048513
9ddfe0ef
00090693
00048713
000a8613
00098593
000c0513
4d0080ef
fff00693
00050d93
00090313
f4d50063
00050463
6140106f
0009a023
00000713
fffff7b7
b0878793
008787b3
0067a023
fffff7b7
b1078793
008787b3
00800613
00000593
000b0513
00e7a023
975fe0ef
040017b7
85078693
fffff7b7
b7878593
b1078793
008787b3
0007a703
0e06a803
fc058793
00070613
000b0693
008785b3
000c0513
000800e7
fffff7b7
b0878793
008787b3
00100693
0007a303
00000713
00d51a63
fffff7b7
fc078793
00878733
b7874703
fffff7b7
fc078793
008787b3
00e78733
b9074703
00071463
47d0106f
00300713
012c8cb3
00ed9463
52c0106f
fffa0a13
fffff7b7
afc78793
008787b3
0007a783
04079663
fffff7b7
af878793
008787b3
0007a783
00498993
02078a63
fffff7b7
af078793
008787b3
0007a783
40f98933
fffff7b7
af478793
008787b3
0007a783
40295713
00f76463
6700106f
004ba703
00000913
00e04463
4f00106f
e20a18e3
fffff7b7
ae878793
008787b3
0007ab03
fffff7b7
afc78793
008787b3
0007a783
06079a63
fffff7b7
af878793
008787b3
0007a783
0009a023
02078c63
fffff7b7
af078793
008787b3
0007a783
40f985b3
fffff7b7
af478793
008787b3
0007a783
4025d713
00170713
00f77463
51d0106f
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
fffff7b7
aec78793
23d0006f
000c0513
6e1070ef
00052783
fffff5b7
af858593
008585b3
00f5a023
fffff7b7
af478793
000016b7
008787b3
fff48713
36c68613
0007a023
02e67263
fffff7b7
c9378713
00e487b3
fffff737
af470713
00870733
00f72023
36d68493
fffff737
aec70713
00870733
00072023
fffff737
af070713
00870733
00072023
fffff737
fffff7b7
b0870713
c9078693
00870733
00072023
fc068713
fffff6b7
00000913
afc68693
780a6993
00000793
00000a13
00870ab3
00023f37
00090713
008686b3
00048913
0166a023
04e00e13
000c0b13
744f0f13
000a0c13
00070493
00098a13
00078993
000ba683
0006c583
fd558713
0ff77713
00ee6a63
00271713
01e70733
00072703
00070067
fffff7b7
af878793
008787b3
0007a783
0007c703
04b71663
200a7713
04070263
fffff7b7
b0878793
008787b3
d7fa7a13
0097a023
00ba8023
fff90913
001a8a93
004ba703
001c8c93
fff70713
00eba223
30e05c63
00168693
00dba023
f80910e3
fffff737
afc70713
00870733
00098793
00048913
000a0993
000c0a13
000b0c13
00072b03
0a048a63
eff9f993
0ac0006f
013c0733
fc0716e3
e7fa7a13
00000993
00000c13
f91ff06f
00100713
faec1ae3
00200c13
f81ff06f
080a7713
fa0702e3
f7fa7a13
f71ff06f
120c16e3
00049a63
700a7713
70000513
00a71463
7440106f
00100713
00e98663
00400713
f6e99ae3
00198993
0ff9f993
f3dff06f
0e0994e3
58049ce3
700a7713
70000513
00a71463
7040106f
fffff737
afc70713
00870733
00098793
000a0993
000c0a13
000b0c13
00072b03
00048913
fffa0e93
00100713
01d76463
2c90106f
fff78713
00600593
66e5f2e3
1009f713
04070063
4009f713
00070463
2dd0106f
fffac583
06500713
fffa8493
fffc8a13
00e58663
04500713
72e59ae3
000b8613
000c0513
19d0c0ef
000a0c93
00048a93
0109f713
a4071663
000a8023
6009f713
40000613
fffff7b7
00c71463
39c0106f
af078793
008787b3
0007a783
00078463
2600106f
fffff7b7
b1078793
008787b3
0007a783
0029f713
0019f993
00478493
600708e3
fffff937
c5090793
00878633
b2090793
00878533
00000693
000c0593
2910b0ef
fc090793
00878733
b6072503
b6472583
b6872603
b6c72683
00099463
1b00106f
00000a13
00000913
fffff7b7
b1078793
008787b3
0007a783
0007a703
01472023
01272223
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
fffff7b7
b1078793
008787b3
000b4703
0097a023
fffff7b7
fc078793
008786b3
b6e6ae23
001b0b13
00070463
fedfe06f
864ff06f
00200793
daf99ae3
00300993
d81ff06f
500a7713
40000793
00f70863
400a7713
d8070ce3
e40484e3
200a7713
02071c63
fffff7b7
b0878793
008787b3
0007a783
fffff737
af070713
40f487b3
00870733
00f72023
fffff7b7
aec78793
008787b3
0157a023
87fa7a13
180a6a13
00000493
d1dff06f
00700793
d4f990e3
00800993
d0dff06f
00600793
d2f998e3
00700993
cfdff06f
100a7713
d40708e3
fffff7b7
af478793
008787b3
0007a783
f7fa7a13
00148493
360794e3
fff90913
cddff06f
000b8593
000b0513
0c10c0ef
000237b7
04e00e13
74478f13
ce0510e3
c4091ce3
cd9ff06f
fffff7b7
af878793
000016b7
008787b3
fff48713
36c68613
0007a023
02e67263
fffff7b7
fffff737
c9378993
af870713
013487b3
00870733
00f72023
36d68493
fffff6b7
b0868693
fffff737
008686b3
c5070793
0006a023
47f70693
00024737
00001937
9b870993
fffff737
d8090a93
b0c70713
015a6ab3
00870733
00878a33
000b0813
000a0b13
00048a13
00072483
000247b7
88078793
80090913
000ba603
04d00513
00064583
fd558713
0ff77713
04e56463
00271713
00f70733
00072703
00070067
00a00713
02975863
00dafab3
00bb0023
001b0b13
004ba703
fff70713
00eba223
16e05663
00160613
00cba023
fffa0a13
fa0a14e3
fffff7b7
b0c78793
008787b3
0097a023
100af713
000b0a13
00080b13
02070663
fffff7b7
c5078793
00878733
01477463
0840106f
fffff7b7
c5078793
00878733
00ea1463
e41fe06f
010af713
4c071463
fffff7b7
c5078793
00878933
fffff7b7
b0c78793
008787b3
0007a683
fffff7b7
b0478793
008787b3
0007a783
00000613
00090593
000c0513
000a0023
000780e7
fffff7b7
b1078793
008787b3
0007a783
020af713
00478993
42071863
008af713
680714e3
004af713
00071463
4900106f
fffff7b7
b1078793
008787b3
0007a783
0007a703
00a71023
4080006f
00149493
009984b3
00049483
00dafab3
eedff06f
600af713
20000513
f0a714e3
dffafa93
500aea93
01000493
ed1ff06f
080af713
ee0708e3
f7fafa93
ec1ff06f
00149493
009984b3
00049483
00800713
ea9744e3
ed1ff06f
012af733
ea0700e3
00049663
200aea93
00800493
400af713
180706e3
a7fafa93
e85ff06f
fffff737
afc70713
00870733
00f72023
fffff7b7
b0c78793
008787b3
000b8593
000c0513
0107a023
62c0c0ef
fffff7b7
47f78693
b0c78793
008787b3
0007a803
fffff7b7
afc78793
008787b3
0007a783
e40508e3
e55ff06f
00049463
00100493
fffff6b7
b0868693
010a7793
008686b3
001a7713
00f6a023
3a070863
00078463
0980106f
fffff7b7
b1078793
008787b3
0007a783
fffff6b7
afc68693
0007a703
008686b3
00478793
00e6a023
fffff6b7
af068693
008686b3
080a7313
00f6a023
00031463
18c0106f
00071463
e41fe06f
08000513
83dfd0ef
00050913
00051463
db9fe06f
fffff7b7
b1c78793
008787b3
fffff6b7
0007a783
afc68693
008686b3
0006a683
0067d983
0047d703
00a6a023
38e9f6e3
0007a503
fffff7b7
b1c78793
008787b3
0007a783
00299713
00198993
01379323
fffff7b7
afc78793
008787b3
0007a783
00e50533
fffff737
00f52023
fffff7b7
af478793
008787b3
af870713
0127a023
00870733
02000793
00f72023
fffff737
b8870993
c9070793
fc070713
00870a33
fc098713
008709b3
fffff737
fc078793
b1070713
008787b3
00870733
00f72023
000b8793
00000a93
000b0b93
00078b13
6e0070ef
59550ee3
000b2783
004b2703
015a06b3
0007c603
fff70713
00178793
00fb2023
c8c68823
00eb2223
00300793
001a8a93
00fd9863
b88a2783
00400713
00e78a63
00800613
00000593
00098513
ee5fd0ef
fffff7b7
b1078793
008787b3
0007a603
00098713
000a8693
00090593
000c0513
1cd070ef
fff00793
00050d93
52f500e3
1c0510e3
fffff7b7
b0878793
008787b3
0007a783
00079463
00092023
015c8cb3
fff48493
fffff7b7
b0878793
008787b3
0007a783
04079463
fffff7b7
afc78793
008787b3
0007a783
02078863
fffff7b7
af478793
008787b3
fffff737
0007a783
af870713
00870733
00072703
40f90ab3
402ad793
18e7f0e3
00490913
004b2783
00000a93
14f056e3
ee049ae3
000b0793
000b8b13
00078b93
fffff7b7
afc78793
008787b3
0007a783
02078a63
fffff7b7
af478793
008787b3
0007a783
40f905b3
fffff7b7
af878793
008787b3
0007a783
4025d713
00f77463
2b40106f
fffff7b7
b0878793
008787b3
0007a783
fffff737
b1870713
0017ba93
fffff7b7
b1878793
008787b3
0007a783
00870733
015787b3
00f72023
fffff7b7
af078793
008787b3
0007a783
fffff737
b1070713
00870733
00f72023
aa1fe06f
fffff7b7
b1078793
008787b3
0007a783
0007a703
00a72023
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
fffff7b7
b1078793
008787b3
0137a023
fffff7b7
c5078793
00878733
fffff7b7
b0878793
008787b3
0007a783
40ea04b3
000b4703
00f484b3
fffff7b7
fc078793
008786b3
b6e6ae23
009c8cb3
001b0b13
00070463
8b1fe06f
929fe06f
ffd98713
0fd77713
e6071a63
f00ff06f
00200793
eefc1463
00300c13
e34ff06f
fffff7b7
b0878793
008787b3
0007a783
480798e3
fffff7b7
b1078793
008787b3
0007a783
080a7313
0007aa83
00478993
62030063
000a9463
8cdfe06f
00048513
ca8fd0ef
00050793
00051463
a25fe06f
fffff737
b1c70713
00870733
00072683
00aaa023
0066d903
0046d703
0006a503
06e96463
fffff6b7
b1068693
008686b3
00f6a023
000106b7
ff668693
00e6f463
9f9fe06f
00870713
01071a13
010a5a13
002a1593
6dd080ef
00051463
9ddfe06f
fffff7b7
b1c78793
008787b3
0007a683
fffff7b7
b1078793
008787b3
0007a783
00a6a023
01469223
fffff6b7
b1c68693
008686b3
0006a683
00291713
00e50733
00190913
01269323
01572023
00048693
000b8713
00100613
00078593
000c0513
18c0c0ef
00050913
00051463
2900106f
54957a63
000aa503
00090593
655080ef
54050263
00aaa023
53c0006f
fffff7b7
afc78793
008787b3
0007a783
280790e3
fffff7b7
b1078793
008787b3
0007a783
fffff737
b1070713
0007aa83
00870733
00478793
080a7313
00f72023
4e0308e3
000a9463
f80fe06f
02000513
b5cfd0ef
00050913
00051463
8d9fe06f
fffff7b7
b1c78793
008787b3
0007a783
00aaa023
0067d983
0047d703
0007a503
70e9f263
fffff7b7
b1c78793
008787b3
0007a783
00299713
00e50533
00198993
01379323
01552023
02000a13
000ba703
fffff7b7
fc078793
00074683
008787b3
00d786b3
b906c683
00069463
efcfe06f
fffff7b7
b0878793
008787b3
0167a023
00090993
000a8b13
000a0a93
0400006f
41378a33
00078913
095a7863
fff48493
2a048663
004ba783
04f05863
000ba703
fffff6b7
fc068693
00074783
008686b3
00f687b3
b907c783
28078263
004ba783
00170693
00dba023
fff78793
00fba223
00074703
00190793
00e90023
fa0b12e3
00078913
fa9ff06f
000b8593
000c0513
7910b0ef
fa0504e3
fffff7b7
b0878793
008787b3
000a8a13
000b0a93
0007ab03
25391263
f8cfe06f
001a9a93
00098513
000a8593
4b1080ef
00050993
00051463
f94fe06f
01450933
00ab2023
f51ff06f
440910e3
fffff7b7
b1078793
008787b3
0007a783
080a7313
0007a983
00478913
24030ee3
00099463
df0fe06f
02000513
9ccfd0ef
00050793
00051463
f48fe06f
fffff737
b1c70713
00870733
00072683
00a9a023
0066da03
0046d703
0006a503
38ea7063
002a1713
00e50533
fffff737
b1c70713
00870733
00072703
001a0a13
01352023
01471323
02000a13
000ba703
00074683
00dd06b3
0006c683
0086f693
02069ce3
fffff6b7
b1068693
008686b3
00078613
0126a023
004ba683
00170593
00bba023
fff68693
00dba223
00074703
00160a93
00e60023
00098663
40fa8933
63497863
fff48493
04048e63
004ba703
02e05263
000ba703
00074683
00dd06b3
0006c683
0086f693
02069e63
000a8613
fa9ff06f
fffff737
b0870713
00870733
000b8593
000c0513
00f72023
6150b0ef
fffff7b7
b0878793
008787b3
0007a783
fa050ae3
fffff737
b1070713
00870733
00072903
40fa84b3
00148593
009c8cb3
000a8793
00078023
00098463
6345e263
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
fffff7b7
b1078793
008787b3
0127a023
d54fe06f
fffff737
afc70713
00098793
00870733
000a0993
00048913
000c0a13
eff9f993
000b0c13
00072b03
a78ff06f
fffff7b7
af478793
008787b3
0007a783
fffff737
af470713
fff78793
00870733
00f72023
958ff06f
fffff7b7
b0878793
008787b3
000a8a13
000b0a93
0007ab03
413904b3
01391463
bfcfe06f
00090023
000a8e63
00148593
0145fa63
000aa503
261080ef
00050463
00aaa023
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
009c8cb3
c90fe06f
fffff737
af870713
00870733
00072703
c7fafa93
00070e63
fffff5b7
af858593
fff70713
008585b3
00e5a023
001a0a13
fffff737
b0870713
00870733
00072703
fffff5b7
b0858593
00170713
008585b3
00e5a023
cb4ff06f
00200713
58f774e3
00300713
98e78a63
ffc78613
0ff67493
fff4ca13
014a8a33
fffac583
000b8613
fffa8a93
000c0513
3450b0ef
ff5a16e3
fffc8813
40980cb3
960ff06f
fffff7b7
c5078793
00000613
008785b3
000c0513
1790a0ef
00050a13
00058913
a0099e63
00050613
00058693
6e8190ef
fffff7b7
b1078793
008787b3
0007a783
0007a983
4e0518e3
000a0513
00090593
5811c0ef
00a9a023
a00ff06f
000b8713
00048693
00100613
000a8593
000c0513
4390b0ef
00050913
00051463
bdcfe06f
fffff7b7
b1878793
008787b3
0007a783
fffff737
b1870713
00178793
00870733
00f72023
fffff7b7
b1078793
008787b3
012c8cb3
0137a023
b38fe06f
000b8613
000c0513
26d0b0ef
ffeac583
ffea8493
ffec8a13
8b8ff06f
fffff6b7
b1068693
008686b3
00f6a023
000106b7
ff668693
00e6f463
ba0fe06f
00870713
01071a93
010ada93
002a9593
085080ef
00051463
b84fe06f
fffff7b7
b1c78793
008787b3
0007a683
fffff7b7
b1078793
008787b3
0007a783
00a6a023
01569223
c21ff06f
fffff6b7
b0868693
008686b3
00f6a023
000106b7
ff668693
00e6f463
b38fe06f
fffff7b7
b1c78793
008787b3
0007a783
00870713
01071713
0007a503
fffff7b7
01075713
b1078793
008787b3
00271593
00e7a023
7f8080ef
00051463
af8fe06f
fffff7b7
fffff737
b1c78793
b1070713
008787b3
00870733
0007a783
00072703
00a7a023
00e79223
fffff7b7
b0878793
008787b3
0007a783
c18fe06f
ffe00793
2af51e63
004b2783
daf04863
000b0593
000c0513
2450b0ef
ea050663
000b0793
000b8b13
00078b93
ea0a8663
a4cfe06f
fffff7b7
af478793
008787b3
0007a503
00371593
768080ef
fffff737
af470713
00870733
00a72023
00051463
a40fe06f
fffff737
afc70713
00870733
fffff7b7
00072703
af878793
008787b3
0007a783
00a72023
fffff737
af870713
00179793
00870733
01550933
00f72023
e18ff06f
000106b7
ff668693
00e6f463
a08fe06f
fffff7b7
b1c78793
008787b3
0007aa83
00870713
01071a13
000aa503
010a5a13
002a1593
6d8080ef
00051463
9d8fe06f
00aaa023
014a9223
c34ff06f
000106b7
ff668693
00e6f463
9bcfe06f
00870713
01071a13
010a5a13
002a1593
6a0080ef
00051463
9a0fe06f
fffff7b7
b1c78793
008787b3
0007a783
00a7a023
01479223
8bdff06f
fffff7b7
b4078793
008787b3
0007a683
00400713
00e68463
ac1fe06f
ac1fe06f
ffe00713
26e518e3
004ba703
00e05463
949fe06f
000b8593
000c0513
0e90b0ef
00051463
b05fe06f
fffff7b7
ae878793
008787b3
0007ab03
00091463
b01fe06f
8e4fe06f
000106b7
ff668693
00e6f463
910fe06f
fffff7b7
b1c78793
008787b3
0007aa83
00870713
01071a13
000aa503
010a5a13
002a1593
5e0080ef
00051463
8e0fe06f
00aaa023
014a9223
82dfe06f
fffff7b7
b1078793
008787b3
0007a783
0007a703
00a70023
d90ff06f
fffff7b7
b1078793
008787b3
0007a783
0007a703
00a72023
00b72223
00c72423
00d72623
e55fe06f
001a1a13
00078513
000a0593
578080ef
00050793
00051463
85cfe06f
01250ab3
00a9a023
9b1ff06f
fffff7b7
aec78793
008787b3
0007aa83
00000613
00a00693
001a8593
000c0513
7090a0ef
fffff7b7
af078793
008787b3
0007a783
40f50633
fb340713
00eae463
fb240a93
000255b7
e8c58593
000a8513
63d080ef
d51fe06f
0009a503
500080ef
9c050ce3
00a9a023
9d1ff06f
00300793
015c8cb3
b8f51c63
b88a2783
00400713
b8e79663
b8cff06f
fffff7b7
af078793
008787b3
0007a503
fffff7b7
af478793
008787b3
0007a783
00379593
4b0080ef
fffff737
af070713
00870733
00a72023
00051463
f89fd06f
fffff737
af870713
00870733
fffff7b7
00072703
af478793
008787b3
0007a783
00a72023
fffff737
af470713
00179793
00870733
012509b3
00f72023
919fe06f
000b0c93
f21fd06f
fffa4583
000b8613
000c0513
fffa0a13
5e00b0ef
f6dfe06f
b0878793
008787b3
0007a783
41278633
f12790e3
c69fe06f
fffff7b7
b7c78993
b1078793
008787b3
0007a783
fffff737
aec70713
00870733
00f72023
fffff7b7
af478793
008787b3
0007a023
fffff7b7
af078793
008787b3
0007a023
fffff7b7
af878793
008787b3
0007a023
fc098793
008789b3
e78fe06f
00100593
889ff06f
000ba683
fffff7b7
fc078793
0006c703
008787b3
00e78733
b9074703
00071463
d19fd06f
004ba703
00168693
00dba023
fff70713
00eba223
00100693
04d48263
04e05463
000ba783
fffff6b7
fc068693
0007c703
008686b3
00e68733
b9074703
02070063
004ba703
00178793
00190913
fff70713
00eba223
00fba023
fd2492e3
012c8cb3
d95fd06f
000b8593
000c0513
5d00b0ef
fa0508e3
012c8cb3
d7dfd06f
fffff737
b0870713
00870733
00072023
fffff737
fffff7b7
afc70713
00870733
b3c78793
00072023
00000a13
00878ab3
fa1fd06f
00000913
0240006f
00e686b3
00dba023
000b8593
000c0513
00e90933
40e484b3
56c0b0ef
2e051c63
004ba703
000ba683
fc974ce3
40970733
009686b3
00990933
00eba223
00dba023
012c8cb3
cf9fd06f
fffff7b7
b1078793
008787b3
0007a783
fffff737
af070713
00870733
00f72023
fffff7b7
af878793
008787b3
0007a023
fffff7b7
af478793
008787b3
0007a023
fffff7b7
afc78793
008787b3
0007a023
00000913
804ff06f
002b4683
008a6a13
002b0b13
b65fd06f
002b4683
002a6a13
002b0b13
b55fd06f
00098793
00000a13
00000993
e04ff06f
ffe00693
00d51463
858fe06f
000aa503
fffff7b7
aec78793
008787b3
0137a023
2ad030ef
fffff7b7
aec78793
008787b3
0007a703
62051663
00300793
013c8cb3
00fd8463
fc1fd06f
fffff7b7
af478793
008787b3
0007a783
b887a703
00400793
00f71463
fa5fd06f
fff90913
f9dfd06f
ff010113
fffff737
00f10793
b1c70713
ff07f793
00870733
00f72023
0007a023
0007a223
a9cfe06f
87fa7a13
00100993
819fe06f
87fa7a13
00100c13
80dfe06f
fffff7b7
afc78793
008787b3
0007a903
fffff7b7
af878793
008787b3
0007a023
fffff7b7
af478793
008787b3
0007a023
fffff7b7
afc78793
008787b3
0007a023
ee1fe06f
000a8913
00000a13
00000a93
b70ff06f
fffff7b7
b1078793
008787b3
0137a023
fffff7b7
b0878793
008787b3
0007a023
fffff7b7
afc78793
008787b3
000a0a93
0007a023
00000a13
d89fd06f
fffff7b7
af878793
008787b3
0007a983
fffff7b7
af478793
008787b3
0007a023
fffff7b7
af078793
008787b3
0007a023
fffff7b7
af878793
008787b3
0007a023
b40fe06f
004a7713
1e070e63
fffff7b7
b1078793
008787b3
01969023
00c7a023
acdfd06f
b1878793
008787b3
0007a023
a11fd06f
000ba683
0006c703
00ed0733
00074703
00877713
04071e63
004ba703
00168693
00dba023
fff70713
00eba223
00100693
00100993
02d48e63
04e05063
000ba783
0007c703
00ed0733
00074703
00877713
02071063
004ba703
00178793
00198993
fff70713
00eba223
00fba023
fd3496e3
013c8cb3
a45fd06f
000b8593
000c0513
2800b0ef
fa050ce3
013c8cb3
a2dfd06f
00091463
a8dfd06f
012c8cb3
a1dfd06f
001af713
00070463
f75fe06f
002afa93
000a9463
f69fe06f
fffff7b7
b0478793
008787b3
0007a783
00011737
b0870713
36e78a63
fffff7b7
b0c78793
008787b3
0007a683
00000613
00090593
000c0513
6800a0ef
00050693
00058713
fffff7b7
b1078793
008787b3
0007a783
0007a603
00d62023
00e62223
f1dfe06f
fffff7b7
ae878793
008787b3
0007ab03
00091463
c08fe06f
fffff7b7
c5078793
00878933
00030493
009907b3
fff7c583
fff48493
000b8613
000c0513
0a00b0ef
fe0494e3
bd8fe06f
00000993
d45fd06f
000a2503
00458593
6e1070ef
00051463
dc1fd06f
00aa2023
db9fd06f
000b0593
000c0513
1700b0ef
00051463
d21fd06f
fffff7b7
af878793
008787b3
0007aa03
fffff7b7
af078793
008787b3
000b8913
000b0b93
0007ab03
00098463
959fd06f
d31fd06f
001a7713
0c071263
002a7313
0a030e63
fffff7b7
b1078793
41fcd713
008787b3
0196a023
00e6a223
00c7a023
8bdfd06f
fffff7b7
af878793
008787b3
0007aa03
fffff7b7
aec78793
008787b3
0007a703
fffff7b7
af078793
008787b3
000b8913
000b0b93
0007ab03
00099463
cc1fd06f
fffff7b7
c5078793
008789b3
00070493
009987b3
fff7c583
fff48493
000b8613
000c0513
7950a0ef
fe0494e3
c91fd06f
fffff7b7
afc78793
008787b3
0007a483
0004a503
5d1070ef
00051463
d35fe06f
00a4a023
d2dfe06f
fffff7b7
b1078793
0196a023
008787b3
00c7a023
80dfd06f
fffff7b7
af878793
008787b3
0007a483
00458593
0004a503
58d070ef
00051463
ac8fe06f
00a4a023
ac0fe06f
fffff4b7
c5048793
008784b3
000b8c93
0154e463
ee8fd06f
fffac583
000c8613
fffa8a93
000c0513
6f50a0ef
fe9a96e3
eccfd06f
fffff4b7
c5048793
008784b3
000b8c93
0154e463
eb4fd06f
fffac583
000c8613
fffa8a93
000c0513
6c10a0ef
fe9a96e3
e98fd06f
fffff7b7
aec78793
008787b3
00e7a023
fffff7b7
afc78793
008787b3
0007a503
fffff7b7
b0878793
008787b3
0007a783
00379593
4dd070ef
fffff737
afc70713
00870733
00a72023
00051463
fb4fd06f
fffff737
aec70713
00870733
00072703
fffff7b7
b0878793
00e50ab3
fffff737
af870713
00870733
00072703
008787b3
0007a783
00a72023
fffff737
b0870713
00179793
00870733
00f72023
acdfd06f
fffff737
b1870713
fff00793
00870733
00f72023
e14fd06f
00025537
e3c50513
45c080ef
00a9a023
d14fe06f
fffff4b7
c5048793
008784b3
000b8c93
0154e463
db4fd06f
fffac583
000c8613
fffa8a93
000c0513
5c10a0ef
fe9a96e3
d98fd06f
fffff7b7
b0c78793
008787b3
0007a683
00000613
00090593
000c0513
2a50a0ef
00050693
00058713
c91ff06f
0009a703
00d70463
f7dfd06f
80cfe06f
fffff7b7
b1878793
008787b3
0007a783
00079463
ec8fd06f
00cbd783
0407f793
00079463
d48fd06f
eb4fd06f
fffff7b7
af878793
008787b3
0007aa03
d65ff06f
e1010113
1e112623
1f212023
1d812423
1da12023
00058c13
00060913
00d12a23
1e812423
1e912223
1d312e23
1d412c23
1d512a23
1d612823
1d712623
1d912223
1bb12e23
00050d13
7a5050ef
00052783
00078513
02f12823
9ccfd0ef
02a12623
0e012823
0e012a23
0e012c23
0e012e23
000d0663
038d2783
70078863
00cc1683
00002637
01069793
0107d793
00c7f5b3
02059863
064c2583
00c6e7b3
01079793
ffffe6b7
4107d793
fff68693
00d5f6b3
00fc1623
01079793
06dc2223
0107d793
0087f693
2e068663
010c2683
2e068263
01a7f793
00a00693
2ed78e63
10c10793
00078893
0ef12223
000247b7
9dc78793
00f12c23
000247b7
bf078793
00090b13
00f12423
000b4783
0e012623
0e012423
02012023
02012a23
02012c23
02012e23
04012223
04012423
00012623
00088c93
22078263
000b0413
02500713
30e78463
00144783
00140413
fe079ae3
416404b3
21640263
0ec12703
0e812783
016ca023
00970733
00178793
009ca223
0ee12623
0ef12423
00700713
008c8c93
2cf74c63
00c12703
00044783
00970733
00e12623
1c078263
fff00313
00144483
0c0103a3
00140413
00000993
00000a13
05a00913
00900a93
02a00b93
00030d93
00140413
fe048793
04f96463
01812703
00279793
00e787b3
0007a783
00078067
00000993
fd048693
00044483
00299793
013787b3
00179793
00f689b3
fd048693
00140413
fedaf2e3
fe048793
fcf970e3
14048463
14910623
0c0103a3
00100a93
00100b93
14c10b13
00012823
00000313
02012423
02012223
00012e23
002a7f93
000f8463
002a8a93
084a7913
0ec12783
00091663
415986b3
44d04ee3
0c714703
02070a63
0e812703
0c710693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
2ee6ca63
020f8a63
0e812703
0c810693
00dca023
00278793
00200693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
52e6c0e3
08000713
22e900e3
41730db3
31b040e3
100a7713
0c071ee3
0e812703
017787b3
016ca023
00170713
017ca223
0ef12623
0ee12423
00700693
3ae6ce63
008c8c93
004a7a13
000a0663
415984b3
3c904463
0159d463
000a8993
00c12703
01370733
00e12623
360790e3
01012783
0e012423
00078863
01012583
000d0513
8c5fb0ef
10c10c93
00040b13
000b4783
de0792e3
0ec12783
00078463
2ed0106f
00cc5783
0407f793
00078463
2240206f
1ec12083
1e812403
00c12503
1e412483
1e012903
1dc12983
1d812a03
1d412a83
1d012b03
1cc12b83
1c812c03
1c412c83
1c012d03
1bc12d83
1f010113
00008067
000c0593
000d0513
780020ef
00050463
1d00206f
00cc5783
00a00693
01a7f793
d0d796e3
00ec1783
d007c2e3
01412683
00090613
000c0593
000d0513
480020ef
00a12623
f7dff06f
000d0513
3f1050ef
00452783
00078513
04f12423
e19fc0ef
00050793
000d0513
00078493
04f12223
3cd050ef
00852783
02f12e23
720492e3
00044483
d89ff06f
00044483
020a6a13
d7dff06f
416404b3
d16416e3
00044783
d41ff06f
0e410613
000c0593
000d0513
1b00f0ef
ee051ee3
10c10c93
d15ff06f
008a7793
000d8313
70079ee3
01412783
0b010513
01b12823
00778793
ff87f793
0047a603
0007a583
00878793
00f12a23
1411b0ef
0b012603
0b412683
0b812703
0bc12783
01012303
0f010513
00612823
0ef12e23
0ec12823
0ed12a23
0ee12c23
29d050ef
0ca12623
00200793
01012303
00f51463
2900106f
00100793
00f51463
3e00106f
06100793
00f49463
7650106f
04100793
00f49463
1850106f
fdf4f713
fff00793
02e12423
00f31463
19c0206f
04700793
00f71463
1800206f
0fc12d83
05412023
0f012e03
0f412e83
0f812f03
100a6793
000dd463
6b90106f
04012c23
00078a13
00012823
fbf48793
02500713
00f77463
5fc0106f
00024737
00279793
b4870713
00e787b3
0007a783
00078067
0e410613
000c0593
000d0513
04612623
05f12023
07c0f0ef
100512e3
0ec12783
04c12303
04012f83
10c10c93
ce5ff06f
0e812483
02012683
00100713
016ca023
00178793
00148493
008c8d93
3ad75ae3
00100713
00eca223
0ef12623
0e912423
00700713
769740e3
02c12703
03012683
00148493
00e787b3
00eda223
00dda023
0ef12623
0e912423
00700713
008d8d93
74974ce3
0f012703
0a010593
0b010513
0ae12823
0f412703
00f12e23
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
7f8180ef
02012783
fff78913
01c12783
360500e3
001b0813
00148493
012787b3
010da023
012da223
0ef12623
0e912423
00700713
008d8d93
30974ae3
03812683
0d410713
00148493
00f687b3
00eda023
00dda223
0ef12623
0e912423
00700713
008d8c93
c49758e3
0e410613
000c0593
000d0513
74d0e0ef
7c051a63
0ec12783
10c10c93
c31ff06f
01000693
0e812703
0096c463
6710106f
000246b7
be068d93
01000913
00700a13
00c0006f
ff048493
04995663
01078793
00170713
01bca023
012ca223
0ef12623
0ee12423
008c8c93
fcea5ee3
0e410613
000c0593
000d0513
6e10e0ef
76051463
ff048493
0ec12783
0e812703
10c10c93
fa994ee3
009787b3
00170713
01bca023
009ca223
0ef12623
0ee12423
00700693
bae6d6e3
0e410613
000c0593
000d0513
6990e0ef
72051063
0ec12783
b91ff06f
000d0513
af0fb0ef
8edff06f
01412703
0c0103a3
00100a93
00072783
00470713
00e12a23
14f10623
00100b93
14c10b13
a6dff06f
01412783
0c0103a3
0007ab03
00478913
4c0b00e3
fff00793
00fd9463
04c0106f
000d8613
00000593
000b0513
01b12a23
585050ef
00a12823
01412303
00051463
4ad0106f
01012783
41678bb3
0c714783
fffbca93
41fada93
01212a23
00012823
02012423
02012223
00012e23
015bfab3
00000313
a00784e3
001a8a93
a01ff06f
01412783
0007a983
00478793
2a09d8e3
413009b3
00f12a23
00044483
004a6a13
961ff06f
01412683
020a7793
00468713
300794e3
010a7793
780790e3
040a7793
00078463
5740106f
200a7a13
760a06e3
01412783
00e12a23
00c12703
0007a783
00040b13
00e78023
aa9ff06f
00044483
06c00793
38f48ee3
010a6a13
905ff06f
01412703
ffff87b7
8307c793
0cf11423
00470793
000d8313
00f12a23
00072d83
000257b7
ea478793
02f12a23
00000913
002a6a93
00200793
07800493
00000693
0cd103a3
fff00693
1ed30463
012de6b3
f7fafa13
1c069c63
24031263
18079e63
001afb93
1b010b13
1e0b90e3
0c714783
000b8a93
006bd463
00030a93
00012823
02012423
02012223
00012e23
ee0796e3
8edff06f
00044483
06800793
32f482e3
040a6a13
85dff06f
02b00793
00044483
0cf103a3
84dff06f
00044483
080a6a13
841ff06f
00044483
00140713
01749463
6850106f
fd048693
00070413
00000d93
82dae2e3
00044483
002d9793
01b787b3
00179793
00d78db3
fd048693
00140413
fedaf2e3
801ff06f
00044483
001a6a13
ff0ff06f
0c714783
00044483
fe079263
02000793
0cf103a3
fd8ff06f
000d8313
010a6a13
020a7793
080784e3
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
bffa7a93
00000793
eddff06f
000d8313
010a6a93
020af793
080780e3
01412783
00778b13
ff8b7b13
008b0793
00f12a23
000b2d83
004b2903
00100793
ea9ff06f
00044483
008a6a13
f60ff06f
000d8313
010a6a13
020a7793
7a078e63
01412783
00778b13
ff8b7b13
004b2783
000b2d83
008b0713
00e12a23
00078913
7c07c663
fff00793
000a0a93
02f30463
012de7b3
f7fa7a93
00079e63
02031263
000a8a13
00000313
00000b93
1b010b13
e69ff06f
2c091ce3
00900793
2db7e8e3
030d8d93
1bb107a3
000a8a13
00100b93
1af10b13
e45ff06f
000a0a93
00100693
fcd78ae3
00200693
06d78c63
1b010b13
01d91713
007df793
003ddd93
03078793
01b76db3
00395913
fefb0fa3
012de733
000b0613
fffb0b13
fc071ce3
001af693
06068a63
03000693
06d78663
ffe60613
1b010793
fedb0fa3
40c78bb3
000a8a13
00060b13
dd5ff06f
00100713
00e79463
3410106f
00200713
000a0a93
f8e798e3
03412683
1b010b13
00fdf793
00f687b3
0007c703
004ddd93
01c91793
01b7edb3
00495913
feeb0fa3
012de7b3
fffb0b13
fc079ce3
1b010793
41678bb3
000a8a13
d79ff06f
06500713
9e975ce3
0f012703
0a010593
0b010513
0ae12823
0f412703
04f12023
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
250180ef
04012783
40051463
0e812703
000256b7
ed468693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
2ee6c6e3
0cc12703
02012683
6ad75063
03012703
02c12683
008c8c93
feecac23
0e812703
00d787b3
fedcae23
00170713
0ef12623
0ee12423
00700693
7ee6c663
02012703
fff70493
e8905463
01000693
0e812703
2a96dce3
01000913
00700b93
00c0006f
ff048493
2a9952e3
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
1410e0ef
1c051463
0ec12783
0e812703
10c10c93
fb5ff06f
41598933
df205063
01000613
0e812703
09265463
04812023
01000e13
000c0413
00700d93
00090c13
00030913
00c0006f
ff0c0c13
058e5a63
00812683
01078793
00170713
00dca023
01cca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
00040593
000d0513
0c10e0ef
20051ce3
01000e13
ff0c0c13
0ec12783
0e812703
10c10c93
fb8e4ae3
00090313
000c0913
00040c13
04012403
00812683
012787b3
00170713
00dca023
012ca223
0ef12623
0ee12423
00700693
008c8c93
d2e6d463
0e410613
000c0593
000d0513
04612023
0590e0ef
0e051063
0ec12783
04012303
10c10c93
d00ff06f
01000613
0e812703
07b65463
01000313
00700913
00c0006f
ff0d8d93
05b35a63
00812683
01078793
00170713
00dca023
006ca223
0ef12623
0ee12423
008c8c93
fce95ce3
0e410613
000c0593
000d0513
7f00e0ef
06051c63
01000313
ff0d8d93
0ec12783
0e812703
10c10c93
fbb34ae3
00812683
01b787b3
00170713
00dca023
01bca223
0ef12623
0ee12423
00700693
008c8c93
c6e6d863
0e410613
000c0593
000d0513
79c0e0ef
02051263
0ec12783
10c10c93
c50ff06f
0e410613
000c0593
000d0513
77c0e0ef
c8050a63
01012583
cc058063
000d0513
d5dfa0ef
cb4ff06f
01000613
0e812703
00d64463
5e00106f
00024637
be060d93
05212623
04812823
000d8913
000d0413
000a8d93
01000e13
00098a93
00700293
00048993
05f12023
000c0493
00068d13
000b0c13
00030b13
00c0006f
ff0d0d13
05ae5a63
01078793
00170713
012ca023
01cca223
0ef12623
0ee12423
008c8c93
fce2dee3
0e410613
00048593
00040513
6d80e0ef
7c051c63
01000e13
ff0d0d13
0ec12783
0e812703
10c10c93
00700293
fbae4ae3
000b0313
000d0693
000c0b13
00040d13
00048c13
04012f83
00098493
05012403
000a8993
000d8a93
00090d93
04c12903
00d787b3
00170713
00dca223
01bca023
0ef12623
0ee12423
00700693
008c8c93
aae6d663
0e410613
000c0593
000d0513
04612623
05f12023
64c0e0ef
ec051ae3
0ec12783
04c12303
04012f83
10c10c93
a7cff06f
0e410613
000c0593
000d0513
04612023
6200e0ef
ea0514e3
0ec12783
04012303
10c10c93
ac0ff06f
0cc12603
64c05e63
01c12703
02012683
00070493
38e6ce63
02905663
0e812703
009787b3
016ca023
00170713
009ca223
0ef12623
0ee12423
00700693
008c8c93
56e6c4e3
fff4c713
41f75713
00e4f4b3
01c12703
409704b3
44904663
01c12683
400a7713
00db04b3
0c0714e3
0cc12683
02012703
00e6c663
001a7713
54070ae3
03012703
02c12603
008c8c93
feecac23
0e812703
00c787b3
feccae23
00170713
0ef12623
0ee12423
00700613
00e65463
3b00106f
02012703
00eb0833
40d70633
40980933
01265463
00060913
03205863
0e812703
012787b3
009ca023
00170713
012ca223
0ef12623
0ee12423
00700693
008c8c93
00e6d463
3e80106f
fff94713
41f75713
00e97933
412604b3
9e905863
01000693
0e812703
6296d063
01000913
00700b93
00c0006f
ff048493
60995663
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
4a80e0ef
d20518e3
0ec12783
0e812703
10c10c93
fb5ff06f
001a7613
c4061663
00eca223
0ef12623
0e912423
00700713
ce975a63
0e410613
000c0593
000d0513
4680e0ef
ce0518e3
0ec12783
0e812483
10c10d93
cd0ff06f
cd205663
01000713
65275463
01000b93
00700b13
00c0006f
ff090913
632bda63
00812703
01078793
00148493
00eda023
017da223
0ef12623
0e912423
008d8d93
fc9b5ce3
0e410613
000c0593
000d0513
4000e0ef
c80514e3
0ec12783
0e812483
10c10d93
fb5ff06f
01412703
010a7793
00072d83
00470713
00e12a23
10079463
040a7793
0e078c63
010d9d93
410ddd93
41fdd913
00090793
8207dee3
01b037b3
41200933
40f90933
41b00db3
000a0a93
02d00693
00100793
e84ff06f
01412703
010a7793
00072d83
00470713
00e12a23
0a079263
040a7793
08078a63
010d9d93
010ddd93
00000913
f6cff06f
01412703
010af793
00072d83
00470713
00e12a23
06079063
040af793
04078663
010d9d93
010ddd93
00000913
00100793
e1cff06f
001a7713
00071463
81cff06f
959ff06f
000d8313
f74ff06f
00044483
00f12a23
ebdfe06f
03000793
1af107a3
1af10b13
e18ff06f
200af793
00078463
0ffdfd93
00000913
00100793
dd0ff06f
200a7793
300790e3
00000913
edcff06f
200a7793
2c0798e3
41fdd913
00090793
f44ff06f
03c12783
00044483
00079463
e61fe06f
0007c783
00079463
e55fe06f
400a6a13
e4dfe06f
00c12603
0006a783
00e12a23
41f65693
00c7a023
00d7a223
00040b13
fbdfe06f
01412703
00072783
00470713
00e12a23
0007a603
0047a683
0087a703
00c7a783
904ff06f
00068493
c69044e3
c8dff06f
000d8313
000a0a93
e5cff06f
000257b7
ea478793
000d8313
02f12a23
020a7793
12078863
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
001a7793
00078e63
012de7b3
00078a63
03000793
0cf10423
0c9104a3
002a6a13
bffa7a93
00200793
cccff06f
000257b7
eb878793
000d8313
02f12a23
fa1ff06f
000d8313
da8ff06f
00144483
020a6a13
00140413
d65fe06f
0e410613
000c0593
000d0513
1a80e0ef
a20518e3
0ec12783
10c10c93
ffcff06f
00144483
200a6a13
00140413
d35fe06f
00600793
000d8b93
13b7eee3
00025837
000b8a93
01212a23
ecc80b13
d7dfe06f
01000693
0e812703
4296de63
01000b93
00700d93
00c0006f
ff048493
429bd463
00812683
01078793
00170713
00dca023
017ca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
000c0593
000d0513
1140e0ef
98051ee3
0ec12783
0e812703
10c10c93
fb5ff06f
01412703
010a7793
00072d83
00470713
00e12a23
06079663
040a7793
04078e63
010d9d93
010ddd93
00000913
ec5ff06f
0e410613
000c0593
000d0513
0c00e0ef
940514e3
0ec12783
0e812483
10c10d93
884ff06f
0e410613
000c0593
000d0513
09c0e0ef
920512e3
0ec12783
0e812483
10c10d93
88cff06f
200a7793
08079ae3
00000913
e6dff06f
1b010b13
00000793
00812823
00912e23
000b0413
03312223
000c0b13
000d8493
00090993
03c12d83
400afa13
0ff00b93
00030c13
00078913
0240006f
00a00613
00000693
00048513
00098593
7d8140ef
52098c63
00050493
00058993
00a00613
00000693
00048513
00098593
579140ef
03050513
fea40fa3
00190913
fff40413
fa0a0ee3
000dc683
fad91ae3
fb7908e3
4a099c63
00900793
4a97e863
000c0313
1b010793
000b0c13
00040b13
01c12483
02412983
01012403
03b12e23
03212023
41678bb3
000a8a13
ac4ff06f
0e812703
000256b7
ed468693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
48e6cc63
18061c63
02012683
001a7713
00d76733
00071463
c55fe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
76e6ce63
02012683
00170713
0168a023
00f687b3
00d8a223
0ef12623
0ee12423
00700693
00888c93
00e6c463
bf9fe06f
fa9fe06f
00040d13
00048c13
f80ff06f
0e410613
000c0593
000d0513
6e50d0ef
f6051663
0ec12783
10c10c93
cfcff06f
00812683
009787b3
009ca223
00dca023
00170713
0ef12623
0ee12423
00700693
00e6c463
b9dfe06f
f51fe06f
00040c13
f2cff06f
0f012783
0a010593
0b010513
0af12823
0f412783
0a012023
0a012223
0af12a23
0f812783
0a012423
0a012623
0af12c23
0fc12783
0af12e23
0ad170ef
4e0540e3
0c714783
04700713
38975c63
00025837
e9880b13
00012823
02012423
02012223
00012e23
f7fa7a13
00300a93
00300b93
00000313
00078463
848ff06f
a49fe06f
01412783
00040b13
0007a783
00e12a23
00c12703
00e7a023
b41fe06f
00812703
012787b3
00148493
00eda023
e55fe06f
000b0513
9fdfb0ef
00050b93
fd9fe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
5ee6ce63
e80650e3
ff000693
40c004b3
52d656e3
01000913
00700b93
00c0006f
ff048493
50995ce3
00812683
01078793
00170713
00d8a023
0128a223
0ef12623
0ee12423
00888893
fcebdce3
0e410613
000c0593
000d0513
5590d0ef
de051063
0ec12783
0e812703
10c10893
fb5ff06f
0fc12783
5607c463
0c714783
04700713
3e975ae3
00025837
ea080b13
eddff06f
00812683
009787b3
00170713
00dca023
009ca223
0ef12623
0ee12423
00700693
008c8c93
f4e6d863
0e410613
000c0593
000d0513
4ed0d0ef
d6051a63
0ec12783
10c10c93
f30ff06f
02012703
02412b83
00812e23
00eb0733
05412023
05312623
03512223
02812983
03612423
03c12403
04412a03
04812a83
00700d93
01000913
000c8693
00070b13
080b8663
08099663
fff40413
fffb8b93
0e812703
014787b3
0156a023
00170713
0146a223
0ef12623
0ee12423
00868693
0eedcc63
00044603
409b0cb3
01965463
00060c93
03905663
0e812603
019787b3
0096a023
00160613
0196a223
0ef12623
0ec12423
0ecdc263
00044603
00868693
fffcc513
41f55513
00acf733
40e60cb3
01904c63
00c484b3
f60b9ee3
12098ee3
fff98993
f7dff06f
0e812603
01994863
0580006f
ff0c8c93
05995863
00812703
01078793
00160613
00e6a023
0126a223
0ef12623
0ec12423
00868693
fccddce3
0e410613
000c0593
000d0513
3bd0d0ef
c4051263
ff0c8c93
0ec12783
0e812603
10c10693
fb994ce3
00812703
019787b3
00160613
00e6a023
0196a223
0ef12623
0ec12423
1acdc4e3
00044603
00868693
00c484b3
f65ff06f
0e410613
000c0593
000d0513
3650d0ef
be051663
0ec12783
10c10693
ef1ff06f
0e410613
000c0593
000d0513
3450d0ef
bc051663
00044603
0ec12783
10c10693
f09ff06f
04412783
04812583
00000913
40f40433
00078613
00040513
2f5060ef
001dc583
00a00613
00000693
00b03833
00048513
00098593
010d8db3
2a4140ef
ad1ff06f
00900793
ac97e4e3
b0dff06f
0e410613
000c0593
000d0513
2d50d0ef
b4051e63
0cc12603
0ec12783
10c10c93
b4dff06f
00025837
e9480b13
c6dff06f
00030693
00200613
0b010a93
0d010793
0cc10713
0dc10813
000a8593
000d0513
04612823
04d12623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
0bb12e23
130030ef
02812703
04700793
01c12f03
02012e83
02412e03
04c12683
05012303
00050b13
04f70ae3
04600793
00d50933
10f716e3
00054703
03000793
38f702e3
0a010b93
0cc12783
00f90933
000b8593
000a8513
00612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
0a012023
0a012223
0a012423
0a012623
22c170ef
01c12303
00090693
02050263
0dc12683
0126fe63
03000713
00168793
0cf12e23
00e68023
0dc12683
ff26e8e3
416687b3
02f12023
0cc12703
04700793
00e12e23
02812703
70f70863
02812703
04600793
0af704e3
01c12783
02812603
04100693
fff78b93
0d712623
0ff4f793
00000713
00d61863
00f78793
0ff7f793
00100713
0cf10a23
02b00793
000bda63
01c12783
00100b93
40fb8bb3
02d00793
0cf10aa3
00900793
1377d4e3
0e310a13
000a0913
00a00593
000b8513
e94f90ef
03050793
fef90fa3
000b8513
00a00593
dfcf90ef
000b8a93
06300793
00090d93
00050b93
fff90913
fd57c6e3
03050693
0ff6f693
ffed8793
fed90fa3
2f47f6e3
0d610713
0080006f
0007c683
00d70023
00178793
00170713
ff4798e3
0e510793
0d610713
41b787b3
00f707b3
0d410713
40e787b3
02f12c23
02012703
03812683
00100793
00d70bb3
14e7dee3
02c12783
00fb8bb3
04012783
fffbca93
41fada93
bff7fa13
100a6a13
015bfab3
02012423
02012223
00012e23
05812783
5e078e63
02d00793
0cf103a3
00000313
001a8a93
c8cfe06f
0e410613
000c0593
000d0513
0550d0ef
8c051e63
0ec12783
10c10c93
a80ff06f
00600b93
ec4ff06f
02012703
00eb0833
40d70633
40980933
b1265e63
00060913
b14ff06f
01412783
00e12a23
00c12703
0007a783
00040b13
00e79023
d40fe06f
018d9d93
418ddd93
41fdd913
00090793
c71fe06f
0ffdfd93
00000913
dd8ff06f
0ffdfd93
00000913
bddfe06f
02d00793
0cf103a3
a99ff06f
0e410613
000c0593
000d0513
7bc0d0ef
d08fe06f
0e410613
000c0593
000d0513
7a80d0ef
00050463
82cff06f
0cc12603
0ec12783
0e812703
10c10893
860650e3
9e1ff06f
05800793
03000713
0ce10423
002a6713
0cf104a3
04e12023
06300793
00012823
14c10b13
7c67c663
0fc12d83
fdf4f793
02f12423
04012c23
0f012e03
0f412e83
0f812f03
102a6a13
520dca63
06100793
00f48463
e78fe06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
25c1a0ef
0cc10613
4a4060ef
00058613
00050593
000a8513
6c9190ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
230170ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
691160ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000257b7
ea478793
02f12223
fff30913
06912023
07312423
07912823
07a12a23
07812c23
01c12483
00090c13
04812e23
07412223
06612623
000b0c93
07612e23
00068d13
000e0d93
000e8913
000f0993
0480006f
000b8593
000a8513
02c12023
01f12e23
0bf12c23
0ac12e23
0b612823
0b412a23
0a012023
0a012223
0a012423
0a012623
5e9160ef
fffc0c13
00090f93
00098613
0e050263
400307b7
00048613
000b8593
000a8513
08f12e23
0ba12023
0bb12223
0b212423
0b312623
08012823
08012a23
08012c23
0f8170ef
000a8513
1d1190ef
00050593
00050413
000a8513
0b012a03
0b412983
0b812b03
0bc12903
2c5190ef
0b012683
04c12603
00048593
08d12023
0b412683
000b8513
09412823
08d12223
0b812683
09312a23
09612c23
08d12423
0bc12683
09212e23
08d12623
454180ef
02412783
0a012b03
0a412a03
008786b3
0006c683
0a812f83
0ac12603
05912a23
00dc8023
05812823
fff00793
001c8c93
000b0d13
000a0d93
000f8913
00060993
eefc10e3
06c12303
000b0393
000a0293
3ffe0937
000b8593
000a8513
02612023
00812e23
06012483
05c12403
06412a03
0a712823
06712223
0a512a23
06512023
0bf12c23
05f12e23
0ac12e23
04c12623
0a012023
0a012223
0a012423
0b212623
565160ef
000c8d93
06812983
07012c83
07412d03
07812c03
07c12b03
02012303
44a04663
000b8593
000a8513
46d160ef
02012303
00051863
01c12783
0017f913
42091663
05012783
03000693
00178713
00ed8733
0007c863
001d8d93
fedd8fa3
ffb71ce3
416d87b3
02f12023
a39ff06f
00130693
00200613
941ff06f
00030693
00300613
935ff06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
709190ef
0cc10613
150060ef
00058613
00050593
000a8513
375190ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
6dd160ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
33d160ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000257b7
eb878793
02f12223
cadff06f
02812b03
02012703
02812e23
04012a03
00eb0733
01c12403
04c12983
02412a83
00068c93
00976463
d0dfe06f
00070493
d05fe06f
01c12703
ffd00793
00f74463
02e35463
ffe48493
fdf4f793
02f12423
8e5ff06f
0c714783
00000313
00078463
c94fe06f
e95fd06f
02012783
01c12703
1af74863
04012783
01c12703
0017f793
00070b93
00078663
02c12783
00f70bb3
04012783
4007f793
00078663
01c12783
2ef04863
fffbca93
41fada93
015bfab3
06700493
02012423
02012223
999ff06f
00012823
00078a13
800007b7
01b7cdb3
02d00793
04f12c23
ac1ff06f
04012783
00d50933
0017f793
0a079c63
0dc12683
81dff06f
0e410613
000c0593
000d0513
1d00d0ef
00050463
a55fe06f
00044603
0ec12783
10c10693
00c484b3
da4ff06f
07800793
a2dff06f
0e410613
000c0593
000d0513
19c0d0ef
00050463
a21fe06f
0cc12683
0ec12783
10c10c93
c31fe06f
02d00793
0cf103a3
b20ff06f
00024637
be060d93
ae9fe06f
0c714783
01212a23
02012423
02012223
00012e23
00030a93
00030b93
00000313
00078463
b68fe06f
d69fd06f
00025837
e9c80b13
aecff06f
0a010b93
f0cff06f
0e410613
000c0593
000d0513
11c0d0ef
00050463
9a1fe06f
0cc12483
02012703
0ec12783
10c10c93
40970633
bf1fe06f
04012783
01c12703
0017f793
0067e7b3
2ae05463
22079263
01c12b83
06600493
04012783
4007f793
18079a63
fffbca93
41fada93
015bfab3
ea5ff06f
000246b7
be068d93
9f0fe06f
02012783
02c12703
06700493
00e78bb3
01c12783
fcf042e3
40fb8bb3
001b8b93
fffbca93
41fada93
015bfab3
e69ff06f
fff00793
00f12623
dd9fd06f
00812683
009787b3
00170713
00d8a023
0098a223
0ef12623
0ee12423
00700693
00888893
92e6d263
0e410613
000c0593
000d0513
0400d0ef
00050463
8c5fe06f
0ec12783
0e812703
10c10893
8fcff06f
0d610793
00071863
03000793
0cf10b23
0d710793
1b010713
030b8b93
40e78733
01778023
0dd70793
02f12c23
f3cff06f
05412783
000d8713
0cf12e23
02412783
fffdc683
00f7c603
02d61063
03000593
feb70fa3
0dc12703
fff70793
0cf12e23
fff74683
fed606e3
00168613
03900593
0ff67613
00b68663
fec70fa3
badff06f
02412783
00a7c603
fec70fa3
b9dff06f
00130593
000d0513
00612823
a95f90ef
01012303
00050b13
1a050663
00a12823
819ff06f
000a0a93
c2cfe06f
00030463
e81fd06f
00100313
e79fd06f
00600313
e71fd06f
04012783
0017f793
ea078463
e9cff06f
06700493
03c12603
0ff00713
00064783
14e78a63
01c12683
00000513
00000593
00d7de63
40f686b3
00164783
04078463
00158593
00160613
fee794e3
02c12e23
00d12e23
02b12223
02a12423
02812783
02412703
04412583
00e78533
b99f80ef
01750bb3
fffbca93
41fada93
015bfab3
e54ff06f
00064783
00150513
fbdff06f
02c12783
06600493
00f70bb3
006b8bb3
dd9ff06f
0a010b93
000b8593
000a8513
04612623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
04d12823
0bb12e23
0a012023
0a012223
0a012423
0a012623
6a4160ef
01c12f03
02012e83
02412e03
04c12303
c2050863
05012683
00100793
40d787b3
0cf12623
c20ff06f
00079a63
00100a93
06600493
00100b93
c15ff06f
02c12783
06600493
00178b93
006b8bb3
fffbca93
41fada93
015bfab3
bf5ff06f
00200793
02f12c23
d48ff06f
01412783
0007ad83
00478793
000dd463
fff00d93
00144483
00f12a23
00070413
98dfd06f
02012423
02012223
ee1ff06f
00cc5783
0407e793
00fc1623
b15fd06f
04001737
00050793
9e472503
00060693
00058613
00078593
f98fd06f
00c5d783
0645ae03
00e5d303
01c5a883
0245a803
b8010113
ffd7f793
40000713
46812c23
00f11a23
00058413
07010793
00810593
46912a23
47212823
46112e23
00050913
07c12623
00611b23
03112223
03012623
00f12423
00f12c23
00e12823
00e12e23
02012023
f2cfd0ef
00050493
02055c63
01415783
0407f793
00078863
00c45783
0407e793
00f41623
47c12083
47812403
47012903
00048513
47412483
48010113
00008067
00810593
00090513
d19f80ef
fc0500e3
fff00493
fb9ff06f
fe010113
00812c23
00912a23
01212823
00112e23
01312623
00050913
00058493
00060413
00050663
03852783
14078a63
00c41703
01842683
00877793
00d42423
01071693
0106d693
08078463
01042783
08078063
00002637
00c6f6b3
0ff4f993
0ff4f493
0a068063
00042703
01442683
40f707b3
0ad7de63
00842683
00170613
00c42023
fff68693
00d42423
01370023
01442703
00178793
0cf70863
00c45783
0017f793
00078663
00a00793
0af48e63
01c12083
01812403
01012903
00c12983
00048513
01412483
02010113
00008067
00040593
00090513
134000ef
08051e63
00c41703
00002637
0ff4f993
01071693
0106d693
00c6f6b3
01042783
0ff4f493
f60694e3
06442683
00c76733
ffffe637
fff60613
00c6f6b3
00e41623
00042703
06d42223
01442683
40f707b3
f4d7c6e3
00040593
00090513
bd1f80ef
02051e63
00042703
00842683
00100793
00170613
fff68693
00c42023
00d42423
01370023
01442703
f2f71ce3
00040593
00090513
b99f80ef
f2050ee3
fff00493
f35ff06f
fd1f80ef
eadff06f
04001737
00050793
9e472503
00058613
00078593
e65ff06f
ff010113
00058713
00812423
00912223
00060593
00050413
042594b7
00068613
00070513
00112623
b404a823
f2cf80ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
040017b7
9e47a783
ff010113
00812423
00912223
00112623
00050493
00058413
00078663
0387a703
08070463
00c41703
01071793
00877693
0107d793
08068863
01042683
0a068863
0017f613
02060863
01442603
00042423
00000513
40c00633
00c42c23
02068a63
00c12083
00812403
00412483
01010113
00008067
0027f613
00000593
00061463
01442583
00b42423
00000513
fc069ae3
0807f793
fc0786e3
04076713
00e41623
fff00513
fbdff06f
00078513
e91f80ef
00c41703
01071793
00877693
0107d793
f6069ce3
0107f693
08068263
0047f793
04079463
01042683
00876713
01071793
00e41623
0107d793
f4069ce3
2807f613
20000593
f4b606e3
00040593
00048513
534030ef
00c41703
01042683
01071793
0107d793
f2dff06f
03042583
00058e63
04040793
00f58863
00048513
f99f80ef
00c41703
02042823
01042683
fdb77713
00042223
00d42023
f91ff06f
00900793
00f4a023
04076713
00e41623
fff00513
f01ff06f
fd010113
000257b7
01412c23
0d07aa03
03212023
02112623
148a2903
02812423
02912223
01312e23
01512a23
01612823
01712623
01812423
04090063
00050b13
00058b93
00100a93
fff00993
00492483
fff48413
02044263
00249493
009904b3
040b8463
1044a783
05778063
fff40413
ffc48493
ff3416e3
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
00492783
0044a683
fff78793
04878e63
0004a223
fa0688e3
18892783
008a9733
00492c03
00f777b3
02079263
000680e7
00492703
148a2783
01871463
f92784e3
f80788e3
00078913
f5dff06f
18c92783
0844a583
00f77733
00071c63
000b0513
000680e7
fcdff06f
00892223
fa9ff06f
00058513
000680e7
fb9ff06f
ff010113
00812423
00912223
00050413
042594b7
00058513
00112623
b404a823
5b1120ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
ff010113
00112623
00812423
00912223
01212023
02058063
00058413
00050493
00050663
03852783
0a078c63
00c41783
02079263
00c12083
00812403
00000913
00412483
00090513
00012903
01010113
00008067
00040593
00048513
d4cf80ef
02c42783
00050913
00078a63
01c42583
00048513
000780e7
06054c63
00c45783
0807f793
06079e63
03042583
00058c63
04040793
00f58663
00048513
d41f80ef
02042823
04442583
00058863
00048513
d2df80ef
04042223
badf80ef
00041623
ba9f80ef
00c12083
00812403
00412483
00090513
00012903
01010113
00008067
b75f80ef
00c41783
f40786e3
f69ff06f
00c45783
fff00913
0807f793
f80786e3
01042583
00048513
cd5f80ef
f7dff06f
040017b7
00050593
9e47a503
ee5ff06f
ff010113
00812423
00000793
00000413
40f40433
00912223
00112623
40245493
02048063
ffc40413
00f40433
00042783
fff48493
ffc40413
000780e7
fe0498e3
00c12083
00812403
00412483
01010113
00008067
00862783
32078063
00c5d683
fd010113
02812423
01412c23
01712623
02112623
02912223
03212023
01312e23
01512a23
01612823
01812423
01912223
01a12023
0086f793
00060b93
00050a13
00058413
08078663
0105a783
08078263
0026f793
000ba483
08078c63
02442783
01c42583
80000ab7
00000993
00000913
c00aca93
00098613
000a0513
04090263
00090693
012af463
000a8693
000780e7
26a05a63
008ba783
00a989b3
40a90933
40a787b3
00fba423
20078863
02442783
01c42583
00098613
000a0513
fc0912e3
0004a983
0044a903
00848493
fa9ff06f
00040593
000a0513
ab9ff0ef
3c051663
00c45683
000ba483
0026f793
f60798e3
0016f793
12079e63
00042783
00842703
80000ab7
ffeacb13
00000c13
00000993
fffaca93
00078513
00070c93
10098263
2006f613
24060e63
00070d13
2ee9ec63
4806f713
08070a63
01442603
01042583
00161713
00c70733
40b78933
01f75c93
00ec8cb3
00190793
401cdc93
013787b3
000c8613
00fcf663
00078c93
00078613
4006f693
2e068463
00060593
000a0513
ff5f80ef
00050d13
30050863
01042583
00090613
4fc030ef
00c45783
b7f7f793
0807e793
00f41623
012d0533
412c87b3
01a42823
01942a23
00a42023
00098c93
00f42423
00098d13
000d0613
000c0593
5e8030ef
00842703
00042783
00098913
41970733
01a787b3
00e42423
00f42023
00000993
008ba783
012c0c33
412787b3
00fba423
0a078a63
00042783
00842703
00c45683
00078513
00070c93
f00992e3
0004ac03
0044a983
00848493
ee9ff06f
00000a93
00000513
00000c13
00000993
0e098063
0e050863
000a8793
00098b13
0137f463
00078b13
00042503
01042783
00842903
01442683
00a7f663
00d90933
0f694263
1adb4e63
02442783
01c42583
000c0613
000a0513
000780e7
00050913
06a05a63
412a8ab3
00100513
040a8c63
008ba783
012c0c33
412989b3
412787b3
00fba423
f80796e3
00000513
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00012d03
03010113
00008067
00040593
000a0513
b90f80ef
fa0500e3
00c41783
0407e793
00f41623
fff00513
fa9ff06f
00000513
00008067
0044a983
00048793
00848493
fe098ae3
0007ac03
00098613
00a00593
000c0513
288030ef
14050463
00150513
41850ab3
ef9ff06f
000c0593
00090613
45c030ef
00042783
00040593
000a0513
012787b3
00f42023
b18f80ef
f0050ee3
f89ff06f
01042683
04f6e863
01442903
0529e463
00098513
013b7463
000a8513
00090593
fa1f70ef
00090593
f75f70ef
02442783
01c42583
00050693
000c0613
000a0513
000780e7
00050913
f2a05ee3
412989b3
e25ff06f
00070913
00e9f463
00098913
00078513
00090613
000c0593
3cc030ef
00842703
00042783
41270733
012787b3
00e42423
00f42023
fc0712e3
00040593
000a0513
a78f80ef
ee0516e3
412989b3
dd5ff06f
00098c93
00098d13
d9dff06f
000b0613
000c0593
380030ef
00842703
00042783
000b0913
41670733
016787b3
00e42423
00f42023
e3dff06f
000a0513
7a4040ef
00050d13
d40510e3
01042583
000a0513
fe8f80ef
00c41783
00c00713
00ea2023
f7f7f793
e81ff06f
00198793
00078a93
db9ff06f
00c00713
00c41783
00ea2023
e65ff06f
fff00513
e11ff06f
00000593
61c0e06f
00450693
00000793
01a50513
ffff8837
01c0006f
00179793
00e69023
01079793
00268693
0107d793
02d50e63
0006d703
00177613
00060463
0017e793
00175713
0027f613
010765b3
fc0606e3
00179793
00b69023
01079793
00268693
0107d793
fcd516e3
00008067
01850693
00000713
00250513
01c0006f
00171713
00f69023
01071713
ffe68693
01075713
04d50463
0006d783
01079613
41065613
00179793
00065463
00176713
01079793
0107d793
00277613
0017e593
fc0600e3
00171713
00b69023
01071713
ffe68693
01075713
fcd510e3
00008067
fc010113
03312623
000109b7
02812c23
02912a23
03212823
03412423
03512223
02112e23
00050a13
00060493
00011d23
00011e23
01858913
01c10413
00810a93
fff98993
00095503
000a0593
ffe40413
ffe90913
02050a63
d35f70ef
00245703
00045683
013577b3
00e787b3
01055513
0107d713
00d50533
00e50533
00a41023
00f41123
01055513
fea41f23
fb541ce3
00448613
01e10713
00045783
00240413
00260613
fef61f23
fee418e3
03c12083
03812403
03412483
03012903
02c12983
02812a03
02412a83
04010113
00008067
00055703
00255783
00070663
00008737
00e7e7b3
00f59923
00255703
000087b7
fff78793
02f70463
00650793
01058593
01850513
0007d703
00278793
ffe58593
00e59123
fea798e3
00008067
00650793
01a50513
0007d703
00278793
02071a63
fea79ae3
01258713
00058793
00278793
fe079f23
fef71ce3
0125d783
00008737
fff70713
00e7e7b3
00f59923
00008067
01058713
00058793
00278793
fe079f23
fef71ce3
ffffc7b7
00f59823
ffff87b7
fff7c793
00f59923
00008067
00455783
ff010113
00912223
00112623
00812423
01212023
00050493
0c079c63
00655703
00000413
01071793
4107d793
0a07c463
01a50693
0a000613
02071863
00648793
0080006f
0007d703
00278793
fee79e23
fed79ae3
00049c23
01040413
06c40c63
0064d703
fc070ce3
f0077793
04079063
01848513
00248593
00000793
00050713
00075683
ffe70713
00869613
00c7e7b3
00f71123
0086d793
feb714e3
0064d703
00840413
f0077793
fc0788e3
0a000913
0140006f
00140413
d49ff0ef
00894c63
0064d703
01071713
41075713
00048513
fe0752e3
00c12083
00040513
00812403
00412483
00012903
01010113
00008067
f007f713
00000413
04071063
f6f00913
0140006f
fff40413
c91ff0ef
fd2404e3
0044d783
00048513
fe0796e3
00c12083
00040513
00812403
00412483
00012903
01010113
00008067
00450693
01a50593
00000713
0080006f
0006d783
0087d613
00c76733
00879793
00e69023
01079713
00268693
01075713
fed590e3
0044d783
ff800413
f89ff06f
fe010113
00812c23
00912a23
00112e23
01212823
01312623
00058493
00050413
0a05c463
00f00793
00058613
00450513
01840693
00f00593
0297d463
00050793
0027d703
00278793
fee79f23
fef69ae3
00041c23
ff060613
fec5c2e3
00f4f493
00700793
0297d863
01840713
00240593
00000793
00075683
ffe70713
00869613
00c7e7b3
00f71123
0086d793
fee594e3
ff848493
00048a63
fff48493
00040513
be9ff0ef
fe049ae3
01c12083
01812403
01412483
01012903
00c12983
00000513
02010113
00008067
ff100793
40b00933
08f5de63
01850593
00000993
00450693
00f00613
01845703
00058793
00e9e9b3
ffe7d703
ffe78793
00e79123
fed79ae3
00041223
ff090913
fd264ee3
ff000913
ff100713
40990933
00000793
08e4ce63
00f90933
00700793
0527ca63
02090063
01845783
fff90913
00040513
0017f793
00f9e9b3
addff0ef
fe0914e3
01c12083
01812403
01412483
01012903
01303533
00c12983
02010113
00008067
ff900793
00000993
00450693
faf5dce3
01844783
01a40593
00f9e9b3
00000793
0006d703
00268693
00875613
00c7e7b3
00871713
fef69f23
01071793
0107d793
feb690e3
ff890913
f79ff06f
ff097793
40f007b3
00f90933
00700793
f727d2e3
fb1ff06f
01255783
00008637
fff60613
00f7d793
40f007b3
00f59023
01255683
01050793
00458713
00c6f6b3
00d59123
02c68663
00658713
00059223
ffe50513
0007d683
ffe78793
00270713
fed71f23
fef518e3
00059c23
00008067
01255603
00d67633
00d61e63
01250813
00050693
0006d603
00268693
00061e63
ff069ae3
01a58593
00270713
fe071f23
fee59ce3
00008067
00658713
00059223
ffc50513
0007d683
ffe78793
00270713
fed71f23
fea798e3
00008067
01255783
fb010113
04812423
fff7c793
04112623
01179713
00058413
00071e63
01250693
00050793
0007d703
00278793
08071c63
fed79ae3
01245783
fff7c793
01179713
06070063
00810593
f01ff0ef
02410593
00040513
ef5ff0ef
00815583
02415503
06b50c63
00a10793
02610713
02010613
0007d683
00278793
0a069863
00075683
00270713
0a069263
fef614e3
00000513
04c12083
04812403
05010113
00008067
00040793
0007d703
01240693
00278793
00071a63
f8d788e3
0007d703
00278793
fe070ae3
04c12083
04812403
ffe00513
05010113
00008067
00a15603
02615683
00153513
00a10713
02610793
00151513
fff50513
03c10593
00278793
00270713
00d61e63
f8b784e3
00075603
0007d683
00270713
00278793
fed606e3
f6c6eae3
40a00533
f6dff06f
00100513
f60582e3
fff00513
f5dff06f
fd010113
02812423
03212023
01312e23
01412c23
01512a23
01712623
00078913
00068b93
02112623
02912223
01612823
00050413
00058993
00060a13
00070a93
a85ff0ef
09000793
40ab8bb3
14a7d463
000087b7
ffe78793
2777d263
220a8c63
00492a83
00092683
01a90713
03490793
2ada8063
00270713
fe071f23
fee79ce3
03800793
32fa8263
1357d863
04000793
2afa8863
07100793
32fa9663
00008737
fff70713
000045b7
01400b13
00a00493
000087b7
00a00613
00860693
00169693
00e91a23
00992423
00b91b23
00f91c23
00c92623
00d90733
00f71523
01592023
01640b33
23705e63
000b5783
01495703
08f00693
00e7f633
0356cc63
00b00693
0296c863
00149713
00e40733
01840693
00275783
00078463
00166613
00071123
00270713
fee696e3
000b5783
01495703
fff74713
00e7f7b3
00fb1023
01695783
00c7f733
0c071463
13705263
00445783
22079663
000087b7
00041c23
ffe78793
1377cc63
01741123
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
03010113
00008067
160bd263
f7000793
12fbdc63
00240793
01a40413
00278793
fe079f23
fe879ce3
fb5ff06f
01800793
1afa8263
03500793
20fa9063
000017b7
7ff00713
40000593
00c00b13
00600493
80078793
00600613
ed5ff06f
01495703
000b5603
fff74793
00f677b3
00fb1023
01695783
00e67633
00c7f733
06070a63
02c79263
18099863
00c92783
01895703
00179793
00f407b3
0007d783
00e7f7b3
f0078ee3
03290513
01840613
01c90913
00000793
00055703
00065803
ffe60613
ffe50513
01070733
00f70733
01075793
00e61123
0017f793
fca91ee3
ef7042e3
09000793
00fa8663
00040513
e50ff0ef
00445783
0e079e63
00041c23
ec0bdee3
00041123
ed9ff06f
00041c23
ffff87b7
fff7c793
00f41123
00440793
01840413
00079023
00278793
fe879ce3
eb1ff06f
00240793
01a40413
00278793
fe079f23
fef41ce3
e99ff06f
000b8593
00040513
965ff0ef
00050463
00100993
d60a9ce3
00041c23
00041123
e75ff06f
e40a8ee3
00492a83
00092683
01a90713
03490793
d6da94e3
00892483
00149b13
01640b33
dd7046e3
09000793
ecfa82e3
01845783
00040513
0017f793
00f9e9b3
d28ff0ef
dadff06f
00010737
fff70713
000085b7
00e00b13
00700493
00100793
00600613
d5dff06f
0ff00713
08000593
00800b13
00400493
10000793
00400613
d41ff06f
00040513
ce0ff0ef
000087b7
001b8b93
00041c23
ffe78793
f177c2e3
ee0bcae3
dc9ff06f
e80a08e3
da5ff06f
0ff00713
08000593
00c00b13
00600493
10000793
00600613
cf9ff06f
00010737
fff70713
000085b7
01800b13
00c00493
00100793
00b00613
cd9ff06f
fd010113
03212023
01312e23
00058913
00255983
02112623
02812423
02912223
01412c23
00060493
01712623
01512a23
01612823
01812423
01912223
01a12023
00050b93
e9cff0ef
00295403
00050793
00090513
40f989b3
03448a13
e84ff0ef
40a40433
04e48713
000a0793
00278793
fe079f23
fee79ce3
09344863
004b8b13
00490a93
01ab8c13
00290d13
000a8713
000b0793
0007d603
00075683
00278793
00270713
0ad61a63
ff8796e3
018b8613
01890713
00000693
00075783
00065583
ffe70713
40d787b3
40b787b3
0107d693
00f71123
0016f693
ffe60613
fced1ee3
00100c93
000a0513
bfcff0ef
04c4d783
fff40413
00090513
00fce7b3
04f49623
be4ff0ef
f93454e3
00040693
02812403
02c12083
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00012d03
00048793
00090513
02412483
02012903
00000713
00000613
00000593
03010113
ac9ff06f
00000c93
f8c6e4e3
f4dff06f
fd010113
02812423
02112623
00058413
00410793
01e10713
00278793
fe079f23
fee79ce3
00e55603
000087b7
fff78793
00f65713
40e00733
00e11223
00f67633
06f60063
00e50793
00c11323
00a10713
ffe7d683
ffe78793
00270713
fed71f23
fef518e3
02061263
00011423
00040593
00410513
c4cff0ef
02c12083
02812403
03010113
00008067
00100793
fff00593
00410513
00f11423
e60ff0ef
fd1ff06f
00050793
00e50693
0007d703
00278793
06071c63
fef69ae3
01440713
00040793
00278793
fe079f23
fee79ce3
01240713
00040793
00278793
fe079f23
fef71ce3
01245783
000086b7
fff68693
00d7e7b3
01079793
0107d793
00f41923
00e51683
f606dce3
00040693
0006d603
00268693
f60614e3
fed71ae3
ffff8737
00e7c7b3
00f41923
f55ff06f
01040713
00040793
00278793
fe079f23
fee79ce3
ffffc7b7
00f41823
ffff87b7
fff7c793
00f41923
f29ff06f
01255783
f5010113
0a812423
fff7c793
0a912223
0b212023
09312e23
0a112623
09412c23
09512a23
09612823
09712623
09812423
09912223
09a12023
07b12e23
01179713
00050493
00058993
00060413
00068913
00071e63
01250693
00050793
0007d703
00278793
2e071a63
fed79ae3
0129d783
fff7c793
01179713
00071e63
01298693
00098793
0007d703
00278793
2e071463
fed79ae3
00024a37
d04a0593
00048513
f84ff0ef
2e050663
0124d603
0129d703
000087b7
fff78793
00f67533
00f775b3
0af51663
01248813
00048793
0007d683
00278793
08069863
ff079ae3
000087b7
fff78793
2cf59263
01298693
00098793
0007d583
00278793
48059663
fed79ae3
01040713
00040793
00278793
fe079f23
fee79ce3
ffffc7b7
00f41823
ffff87b7
fff7c793
00f41923
0ac12083
0a812403
0a412483
0a012903
09c12983
09812a03
09412a83
09012b03
08c12b83
08812c03
08412c83
08012d03
07c12d83
0b010113
00008067
000087b7
fff78793
24f58863
00048513
01c10593
df8ff0ef
03810593
00098513
decff0ef
03a15a83
01e15483
2a0a8e63
01512623
00048713
00912423
02010793
03410693
02071263
38d78c63
0007d703
00278793
fe070ae3
01c10513
a64ff0ef
40a487b3
00f12423
03812703
03890a93
000a8793
02e92a23
04e90493
00278793
fe079f23
fef49ce3
03810513
fd1fe0ef
02215b03
000109b7
05010c13
010b1a13
416a0a33
03a10c93
fff98993
06e10d13
05610d93
03c15503
03e15783
00098b93
01051513
00f50533
00aa6a63
000b0593
e1df60ef
01051b93
010bdb93
05410613
01c10593
000b8513
84cff0ef
03c10713
05810793
0007d603
00075683
00278793
00270713
20d61a63
ffa796e3
00000793
06c10693
000c0613
00065703
0006d583
ffe60613
40f70733
40b70733
01075793
00e61123
0017f793
ffe68693
fd961ee3
017a9023
03c10793
0027d703
00278793
fee79f23
ff879ae3
04011823
002a8a93
f5549ae3
00000713
03c10793
05210613
0007d683
00278793
00d76733
fec79ae3
00e035b3
03810793
03490713
00075683
00278793
00270713
fed79f23
fef618e3
00c12783
00812703
000046b7
fff68693
40e78ab3
03810513
00090793
04000713
00da86b3
00000613
e34ff0ef
03815703
01c15783
00040593
03810513
40e787b3
00f037b3
40f007b3
02f11c23
818ff0ef
dd5ff06f
01448713
0004d783
00248493
00240413
fef41f23
fee498e3
db9ff06f
01440713
0009d783
00240413
00298993
fef41f23
fee418e3
d9dff06f
d04a0593
00098513
c8cff0ef
d00516e3
d61ff06f
dc0806e3
01440793
00240413
fe041f23
fef41ce3
d71ff06f
00000813
01298693
00098793
0007d583
00278793
fc059ae3
fed79ae3
000087b7
fff78793
04f50a63
00f65613
0009d783
00298993
18079263
fed99ae3
00f75793
00c7c7b3
00f79793
00f41923
01240713
00040793
00278793
fe079f23
fee79ce3
01245783
00008737
fff70713
00e7e7b3
00f41923
cf9ff06f
01248593
0004d783
00248493
12079e63
feb49ae3
f9dff06f
03c10793
05010c13
0cfc0e63
0007d703
00278793
fe070ae3
03810513
fbdfe0ef
40a007b3
01e15703
00f12623
d25ff06f
dec6fae3
fffb8793
01079513
01055513
00000693
03410613
06c10713
00075783
00065583
ffe70713
40d787b3
40b787b3
0107d693
00f71123
0016f693
ffe60613
fdb71ee3
03c10713
05810793
0007d603
00075683
00278793
00270713
00d61863
ffa796e3
00050b93
d8dff06f
fec6fce3
ffeb8893
01089b93
010bdb93
00000693
03410613
06c10713
00075783
00065583
ffe70713
40d787b3
40b787b3
0107d693
00f71123
0016f693
ffe60613
fdb71ee3
d45ff06f
01440793
00240413
fe041f23
fef41ce3
be9ff06f
01c15683
03815603
01240713
00040793
40c686b3
00d036b3
00f69693
00d41923
00278793
fe079f23
fef71ce3
eadff06f
00000793
e85ff06f
00000613
e69ff06f
00100813
e3dff06f
f7010113
08912223
00050493
01255503
00008737
fff70713
08812423
09212023
07412c23
08112623
07312e23
07512a23
07612823
07712623
07812423
07912223
00e57833
00058913
00060413
00068a13
00e81e63
01248993
00048713
00075603
00270713
1e061463
ff371ae3
01295603
000087b7
fff78793
00f675b3
08f58863
1ef81463
01248993
00048793
0007d703
00278793
26071663
fef99ae3
000245b7
d0458593
00090513
9f0ff0ef
22050463
01295603
000087b7
fff78793
00f675b3
24f58663
0124d503
00f57733
18f71e63
00048793
0007d703
00278793
3c071063
fef99ae3
0004d783
00248493
36079c63
ff349ae3
00f55713
000087b7
fff78793
0cf59063
01290693
0a80006f
01290693
00090713
00075783
00270713
18079e63
fee69ae3
000087b7
fff78793
f4f80ce3
00090793
0007d703
00278793
0e071863
fef69ae3
000245b7
d0458593
00048513
948ff0ef
18050063
0124d503
01295603
000087b7
fff78793
00f57833
00f675b3
0cf80a63
000087b7
fff78793
0ef59663
01290693
00090793
0007d703
00278793
0c071c63
fed79ae3
000087b7
fff78793
00f55713
00080593
01248993
f2f80ce3
00095783
00290913
2a079a63
fed91ae3
00f65793
00e7c7b3
00f79793
00f41923
01240713
00040793
00278793
fe079f23
fee79ce3
01245783
00008737
fff70713
00e7e7b3
00f41923
08c12083
08812403
08412483
08012903
07c12983
07812a03
07412a83
07012b03
06c12b83
06812c03
06412c83
09010113
00008067
0124d503
000087b7
fff78793
00f575b3
00058813
f4f592e3
01248993
e89ff06f
01440713
0004d783
00240413
00248493
fef41f23
fee418e3
f95ff06f
00048513
00c10593
f75fe0ef
02810593
00090513
f69fe0ef
00e15483
02a15983
08049663
01010793
02410693
1ef68063
0007d703
00278793
fe070ae3
00c10513
bf1fe0ef
02a15703
40a004b3
0640006f
01490713
00095783
00290913
00240413
fef41f23
fee918e3
f29ff06f
01040713
00040793
00278793
fe079f23
fee79ce3
ffffc7b7
00f41823
ffff87b7
fff7c793
00f41923
efdff06f
000087b7
fff78793
dcf594e3
01290693
e21ff06f
00098713
00098913
02c10793
04010693
02071263
16d78063
0007d703
00278793
fe070ae3
02810513
b5dfe0ef
02a15703
40a98933
02815783
038a0993
02ea1b23
02fa1a23
04ea0713
00098793
00079023
00278793
fee79ce3
04ca0c13
00000b93
02410a93
01010c93
04610b13
000ad503
ffea8a93
08051c63
04ca5783
000c0713
00fbebb3
ffe75603
ffe70713
00c71123
fee99ae3
020a1c23
fd9a9ae3
034a0713
02810793
04210613
00075683
00278793
00270713
fed79f23
fec798e3
ffffc6b7
012484b3
00268693
000b8593
02810513
000a0793
04000713
00d486b3
00000613
fe1fe0ef
02815703
00c15783
00040593
02810513
40e787b3
00f037b3
40f007b3
02f11423
9c5fe0ef
dddff06f
04410613
02810593
8e5fe0ef
000c0513
00000593
05c10613
00055783
00065703
ffe50513
ffe60613
00f70733
00b70733
01075593
00e51123
0015f593
fd661ee3
f2dff06f
00000713
c91ff06f
00000793
d55ff06f
01440793
00240413
fe041f23
fef41ce3
d75ff06f
01440793
00240413
fe041f23
fef41ce3
d61ff06f
00008837
fff80813
cd1ff06f
00c5a883
e1010113
0005ae83
0045ae03
0085a303
03112e23
04052583
fff00893
1e812423
17112023
00078413
09000893
09000793
1d412c23
1e112623
1e912223
1f212023
1d312e23
1d512a23
1d612823
1d712623
1d812423
1d912223
1da12023
1bb12e23
03d12823
03c12a23
02612c23
17112223
00c12023
00d12423
00e12823
01012a23
00f12623
00050a13
02058463
04452703
00100793
00e797b3
00f5a423
00e5a223
3b1010ef
16412783
040a2023
00f12623
06010913
00090593
03010513
bb4ff0ef
07215783
00008737
fff70713
00e7f5b3
00e59e63
00090713
07210613
00075683
00270713
3c0694e3
fec71ae3
00f7d793
00012703
00f42023
00300793
08f70ae3
01400793
00f12223
3a0716e3
000087b7
fff78793
00f59e63
00090793
07210693
0007d703
00278793
0e0712e3
fed79ae3
09000793
16f12223
07c10713
00090793
07410613
0007d683
00278793
00270713
fed71f23
fec798e3
08e15603
00012c23
01061793
4107d793
5607c863
00024bb7
d04b8d93
014d8c13
00000693
09810793
000c0713
0ac10d13
0080006f
00075683
00278793
fed79f23
00270713
ffa798e3
14060463
000087b7
fff78793
4af60ee3
08c11783
5207dce3
07c10593
000c0513
c2dfe0ef
12050e63
060542e3
08e15783
5c0796e3
08c11783
00000493
16010993
0207c463
118d8413
07c10613
00098693
00060593
00040513
95dff0ef
08c11783
fff48493
fe07d2e3
0d010413
0e810b13
00040713
07c10793
09010613
0007d683
00278793
00270713
fed71f23
fec798e3
00000693
09810793
000c0713
0080006f
00075683
00278793
fed79f23
00270713
ffa798e3
028d8d13
12cd8c93
fffffab7
21cd8d93
00c0006f
014c8c93
014d0d13
00040593
000c0513
b75fe0ef
04a05863
00040593
000c8513
b65fe0ef
02054863
00098693
00040613
00040593
000d0513
8b5ff0ef
09810613
00098693
00060593
000d0513
8a1ff0ef
015484b3
01fad793
015787b3
4017da93
fbbc90e3
09810613
00098693
000c0593
00060513
ae8ff0ef
12410a93
0300006f
07c10793
08e10693
0007d703
ec0712e3
00278793
fed79ae3
00000493
12410a93
16010993
0d010413
0e810b13
00040593
09810513
a1dfe0ef
09810713
00040793
0007d683
00278793
00270713
fed71f23
ff6798e3
00040593
07c10513
0a011823
9f1fe0ef
07c10793
00045703
00240413
00278793
fee79f23
ff6418e3
09810513
00098613
07c10593
08011a23
f99fe0ef
1ac15503
16051a63
09410c13
07e10c93
0b610413
d04b8593
07c10513
a59fe0ef
14050c63
00000713
000c0693
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fd9690e3
0b410713
07c10793
0007d683
00278793
00270713
fed71f23
ff8798e3
0c011623
00000713
0cc10693
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fc8690e3
00000713
0cc10693
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fc8690e3
00000613
000c0693
0cc10713
0006d583
00075783
ffe68693
ffe70713
00b787b3
00c787b3
0107d613
00f69123
00167613
fc871ee3
09810513
00098613
07c10593
e2dfe0ef
1ac15503
fff48493
ea0500e3
01812783
00012683
00300713
00f037b3
40f007b3
00d7f793
02078793
12f10223
00412783
00e69463
009787b3
02a00713
00f12c23
00f75463
00e12c23
00a00713
4ae50463
03050513
02e00713
12a102a3
12e10323
1c07c4e3
12710b13
00000413
00912e23
000b0493
00040b13
01812403
0b410c93
09410d13
07e10d93
0b610c13
00000693
000d0613
00065783
01079593
4105d593
0005d463
0016e693
00179793
01079793
0026f593
0107d793
00058463
0017e793
00169693
00f61023
01069693
ffe60613
0106d693
fdb610e3
000c8693
07c10793
0007d603
00278793
00268693
fec69f23
ffa798e3
0c011623
00000693
0cc10613
00065783
01079593
4105d593
0005d463
0016e693
00179793
01079793
0026f593
0107d793
00058463
0017e793
00169693
00f61023
01069693
ffe60613
0106d693
fd8610e3
00000693
0cc10613
00065783
01079593
4105d593
0005d463
0016e693
00179793
01079793
0026f593
0107d793
00058463
0017e793
00169693
00f61023
01069693
ffe60613
0106d693
fd8610e3
00000593
000d0613
0cc10693
00065503
0006d783
ffe60613
ffe68693
00a787b3
00b787b3
0107d593
00f61123
0015f593
fd869ee3
00098613
07c10593
09810513
c59fe0ef
1ac15603
00148793
001b0b13
03060693
fed78fa3
03644463
00078493
e9dff06f
01161613
000107b7
01165613
fff78793
08c11723
00f12c23
a7dff06f
00048b13
01c12483
00400713
04c75a63
00500713
00e60ae3
ffe7c703
01812683
ffe78613
07f77713
0206c663
02e00793
03800593
03000513
76f70663
78e5d263
fff64703
00a60023
fff60613
07f77713
fe9ff06f
03100713
fee78f23
00148493
000255b7
00048613
ef458593
000b0513
088030ef
07215783
00c12703
16912823
fff7c793
16e12223
01179713
18070863
01012683
12414703
00148793
00f6a023
000a8793
02070a63
02e00693
20d70663
0017c703
00178793
fe071ae3
04500693
00fae663
0140006f
01578863
fff7c703
fff78793
fed71ae3
00078023
000a8793
02000693
02d00613
0007c703
00d70463
00c71663
00178793
ff1ff06f
000a8413
00c0006f
0007c703
00068413
00e40023
00140693
00178793
fe0716e3
00012703
00200793
fff44683
12f70063
00412783
00078713
0097d463
00048713
03000793
02f69663
415407b3
02f75263
03000693
00c0006f
415407b3
00f75a63
ffe44783
fe040fa3
fff40413
fed786e3
00012703
00300793
0ef70663
00812783
040a2223
00978613
01700793
10c7f663
00100713
00400793
00179793
01478693
00070593
00170713
fed678e3
04ba2223
000a0513
304010ef
00050493
080502e3
04aa2023
000a8593
7b1020ef
01412703
00070863
415407b3
00f487b3
00f72023
1ec12083
1e812403
1e012903
1dc12983
1d812a03
1d412a83
1d012b03
1cc12b83
1c812c03
1c412c83
1c012d03
1bc12d83
00048513
1e412483
1f010113
00008067
00090793
07210693
0007d703
00278793
5a071063
fed79ae3
01012703
000027b7
70f78793
00f72023
e99ff06f
03000793
f2f696e3
415407b3
00100713
eef74ae3
f1dff06f
00412783
009784b3
4e04c063
01012783
00812703
0007a783
00f707b3
00f12423
00812783
040a2223
00378613
01700793
eec7eee3
00000593
f15ff06f
00812783
00078713
00f12223
02a00793
f6e7d663
00f12223
f64ff06f
0007c703
e00700e3
0017c703
00178793
fee78fa3
de0708e3
0017c703
00178793
fee78fa3
fe0712e3
dddff06f
03100713
12e102a3
02e00713
12e10323
00148493
2af05a63
03000793
12f103a3
01812783
12810b13
fff78793
00f12c23
b45ff06f
12410a93
000255b7
f6058593
000a8513
000024b7
5cd020ef
70f48493
d41ff06f
0b410c93
000c8713
07c10793
09010613
0007d683
00278793
00270713
fed71f23
fec798e3
000047b7
08e78793
0cf11323
000087b7
fff78793
00f12e23
ffffc7b7
12410a93
0d010413
01000713
0c8d8313
00278793
03412423
03512223
00000493
00040a93
16010993
0aa10b13
02f12023
00030a13
00070413
00098693
09810613
000c8593
000a0513
b11fe0ef
04c10713
09810793
0007d683
00278793
00270713
fed71f23
ffa798e3
01c12783
05e15583
00f5f533
02012783
00f50533
36a05463
09000613
40a60633
000a8713
04c10793
0007d683
00278793
00270713
fed71f23
ff2798e3
06c05663
00f00793
000a8713
02c7de63
08000693
40a686b3
0046d693
00168713
00171713
00ea8733
000a8793
00278793
fe079f23
fef71ce3
08000613
40a60633
00469693
40d60633
00161793
00fd87b3
00075683
2307d783
00f6f7b3
00f71023
01059593
4105d593
1405c463
09810793
000a8713
0007d603
00075683
02d61863
00278793
00270713
fefb16e3
000c8713
09810793
0007d683
00278793
00270713
fed71f23
ffa798e3
008484b3
014a0a13
12cd8793
00145413
ecfa1ee3
0c615783
08e15703
000a8413
02812a03
00e787b3
ffffc737
f7270713
02412a83
00e787b3
0cf11323
07c10713
000c8793
0c810613
0007d683
00278793
00270713
fed71f23
fec798e3
00000713
09810793
0080006f
000c5703
00278793
fee79f23
002c0c13
ffa798e3
028d8b13
00001c37
118d8d93
0100006f
001c5c13
25bb0463
014b0b13
000c8593
000d8513
994fe0ef
22a04a63
000c8593
000b0513
984fe0ef
fca04ce3
00098693
000c8613
000c8593
000b0513
945fe0ef
09810613
00098693
00060593
000b0513
ec1fe0ef
018484b3
fa9ff06f
12710b13
aa0798e3
8a5ff06f
00000793
c40ff06f
00812783
fff78793
cd9ff06f
04c10793
000a8713
0140006f
00278793
05e10693
00270713
ead782e3
0007d603
00075683
fed604e3
0e215783
01c12703
00e7f7b3
3ce78063
0ec10593
000c0513
838fe0ef
10810593
000a8513
82cfe0ef
0ec15703
10a15603
0ee15883
fff74713
01071713
01075713
0ee11623
40c885b3
00060693
06b05e63
02412583
10810693
12010793
0006d503
00268693
00258593
fea59f23
fef698e3
12011e23
10810693
0ec10593
0080006f
0005d703
00268693
fee69f23
00258593
fef698e3
02412783
12011023
0ec10713
13c10513
0007d683
00278793
00270713
fed71f23
fea798e3
10a15683
411605b3
10011223
00068613
32058c63
02d12623
f6f00793
06f5c863
0ec10513
da5fd0ef
02c12683
00050593
12010793
10410713
0ec15503
10815603
3ac50863
00000613
10a10893
00060513
0007d603
00075803
ffe78793
40a60633
41060633
01065513
00c79123
00157513
ffe70713
fd179ee3
00100613
00098793
04000713
10810513
900fe0ef
000a8593
10810513
afdfd0ef
d45ff06f
01012783
12010223
000a8413
0007a023
b29ff06f
000a8793
0e410713
00278793
fe079f23
fee79ce3
d0dff06f
01812783
12410a93
10078263
000255b7
ed858593
000a8513
000024b7
169020ef
70f48493
8ddff06f
0e810b13
c80ff06f
fff64783
03800713
0ef77863
03100793
00148493
fef60fa3
8a5ff06f
00170713
00e60023
899ff06f
07210713
0080006f
8ae90ee3
00095783
00290913
fe078ae3
01012703
000027b7
70f78793
00f72023
8e9ff06f
12410a93
000255b7
ef058593
000a8513
000024b7
0ed020ef
70f48493
861ff06f
1ac15603
12610b13
12710793
fe4ff06f
09810593
07c10513
00f12e23
a09fd0ef
d04b8593
09810513
eb9fd0ef
01c12783
fc051863
01812703
800748e3
ffe7c703
fd270613
00163613
fff64613
00cb0633
00064603
00167613
fe060863
ffe78613
07f77713
fb0ff06f
000255b7
ee458593
000a8513
000024b7
069020ef
70f48493
fdcff06f
00178793
fef60fa3
fbcff06f
0d010413
00040593
07c10513
00004cb7
d8dfd0ef
00000493
0e810b13
0cc10993
0d210a93
ffec8c93
0e815783
0077f793
0c079a63
0b410713
00040793
0007d683
00278793
00270713
fed71f23
ff6798e3
0b410513
0c011623
f94fd0ef
0b410513
f8cfd0ef
00000613
00098693
000b0713
0006d583
00075783
ffe68693
ffe70713
00b787b3
00c787b3
0107d613
00f69123
00167613
fd571ee3
0b615783
0b815703
00378793
0af11b23
02070063
0b410513
f3cfd0ef
0b615783
0b815703
00178793
0af11b23
fe0714e3
0cc15783
02079c63
0b615783
02fce863
00040713
0b410793
0007d683
00278793
00270713
fed71f23
ff3798e3
0e011423
fff48493
fd500793
f2f494e3
07c10593
00040513
889fd0ef
16010993
960ff06f
000a8793
0007d703
00278793
aa071ee3
0e210713
fee798e3
000a8793
0007d703
00278793
c20710e3
0e210713
fee798e3
a99ff06f
10c10713
0f010793
0007d883
00075503
00278793
00270713
04a89863
10610513
fea794e3
0ec15703
10815783
04f70663
000a8793
0e410713
00278793
fe079f23
fee79ce3
a51ff06f
000256b7
000015b7
00025537
ef868693
00000613
b6e58593
f0c50513
2e90a0ef
07156c63
12010793
10410713
c7dff06f
00068713
00069663
10e11783
0c07d663
10a10713
12010793
00075583
10059663
00270713
fee79ae3
10c11523
ca1ff06f
00000613
0ee10893
0007d803
00075503
ffe78793
ffe70713
01050533
00c50633
01065513
00c79123
00157613
fd171ee3
00000613
c59ff06f
02412603
10810713
12010793
00075503
00270713
00260613
fea61f23
fef718e3
12011e23
10810513
0ec10613
10410713
00065803
00260613
00250513
ff051f23
fee618e3
02412603
12011023
0ec10893
13c10513
00065803
00260613
00288893
ff089f23
fea618e3
10011223
ba5ff06f
12010693
10a10893
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fd1690e3
ba9ff06f
00168613
10c11523
b9dff06f
00852703
00c52783
00052603
00452683
fc010113
00010513
01410593
00e12423
00f12623
02112e23
00c12023
00d12223
9acfe0ef
02615783
00000513
fff7c793
01179713
02071063
01410793
02610693
0007d703
00278793
00071c63
fed79ae3
00200513
03c12083
04010113
00008067
00100513
ff1ff06f
0f050513
00008067
04001537
94050513
00008067
04001537
94050513
00008067
ff010113
00112623
00812423
00912223
02060c63
000255b7
f6c58593
00060513
00060413
880f70ef
000254b7
02051263
f6848513
00c12083
00812403
00412483
01010113
00008067
000254b7
fe5ff06f
f6848593
00040513
84cf70ef
fc050ae3
000255b7
e3c58593
00040513
838f70ef
fc0500e3
00000513
fbdff06f
040017b7
9787c503
00008067
ff010113
00112623
00812423
00912223
02058c63
00058413
000255b7
f6c58593
00040513
ff9f60ef
000254b7
02051263
f6848513
00c12083
00812403
00412483
01010113
00008067
000254b7
fe5ff06f
f6848593
00040513
fc5f60ef
fc050ae3
000255b7
e3c58593
00040513
fb1f60ef
fc0500e3
00000513
fbdff06f
ff010113
00058713
00812423
00912223
00060593
00050413
042594b7
00068613
00070513
00112623
b404a823
3a50f0ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
00c5d783
f8010113
06812c23
06112e23
06912a23
07212823
07312623
07412423
0027f713
00058413
02070c63
04358793
00f5a023
00f5a823
00100793
00f5aa23
07c12083
07812403
07412483
07012903
06c12983
06812a03
08010113
00008067
00e59583
00050493
0805cc63
00810613
3a10a0ef
08054463
00c12783
0000f937
000019b7
00f97933
ffffe7b7
00f90933
00193913
40000a13
80098993
000a0593
00048513
f05f50ef
00c41783
06050e63
00001737
52c70713
02e4ae23
0807e793
00f41623
00a42023
00a42823
01442a23
08091863
0137e7b3
07c12083
00f41623
07812403
07412483
07012903
06c12983
06812a03
08010113
00008067
00c45783
0807f793
00000913
04078663
04000a13
000a0593
00048513
e91f50ef
00c41783
00000993
f80516e3
2007f713
f0071ae3
ffc7f793
0027e793
04340713
00f41623
00100793
00e42023
00e42823
00f42a23
ef1ff06f
40000a13
00000993
f41ff06f
00e41583
00048513
73c0b0ef
00051663
00c41783
f61ff06f
00c45783
ffc7f793
0017e793
01079793
4107d793
f49ff06f
f9010113
06812423
00058413
00e59583
06912223
07212023
06112623
00060493
00068913
0405ca63
00810613
2550a0ef
04054463
00c12703
0000f7b7
06c12083
00e7f7b3
ffffe737
00e787b3
06812403
0017b793
00f92023
40000713
00e4a023
00001537
06412483
06012903
80050513
07010113
00008067
00c45783
0807f793
02078863
06c12083
06812403
00000793
00f92023
04000713
00e4a023
06012903
06412483
00000513
07010113
00008067
06c12083
06812403
00000793
00f92023
40000713
00e4a023
06012903
06412483
00000513
07010113
00008067
ff010113
00812423
00912223
040017b7
00112623
9347a783
00050413
00070493
02060263
000780e7
fff00793
02f50a63
00c12083
00812403
00412483
01010113
00008067
00025637
00100693
e3c60613
00000593
000780e7
fff00793
fcf51ae3
0004a023
08a00793
00c12083
00f42023
00812403
00412483
01010113
00008067
ff010113
04001737
00812423
00912223
00112623
9e472483
04001737
93472803
00068413
02058c63
00060693
00040713
00058613
00050593
00048513
000800e7
fff00793
02f50c63
00c12083
00812403
00412483
01010113
00008067
00025637
00068713
e3c60613
00100693
00048513
000800e7
fff00793
fcf518e3
00042023
00c12083
00812403
08a00793
00f4a023
00412483
01010113
00008067
040017b7
9347a783
00078067
02058063
04060263
04068863
00064783
00f5a023
00064503
00a03533
00008067
ff010113
00c10593
02060463
02068a63
00064783
00f5a023
00064503
00a03533
01010113
00008067
00000513
00008067
00000513
fedff06f
ffe00513
00008067
ffe00513
fddff06f
00357793
0ff5f693
02078a63
fff60793
02060e63
fff00613
0180006f
00150513
00357713
00070e63
fff78793
02c78063
00054703
fed714e3
00008067
00060793
00300713
02f76663
00079663
00000513
00008067
00f507b3
00c0006f
00150513
fea786e3
00054703
fed71ae3
00008067
0ff5f593
00859713
00b76733
01071893
feff0837
808085b7
00e8e8b3
eff80813
08058593
00300313
00052703
00e8c733
01070633
fff74713
00e67733
00b77733
fa0712e3
ffc78793
00450513
fcf36ee3
f8079ae3
f89ff06f
00b547b3
0037f793
00c508b3
06079663
00300793
06c7f263
00357793
00050713
0c079a63
ffc8f613
40e606b3
02000793
02000293
06d7c263
00058693
00070793
02c77863
0006a803
00478793
00468693
ff07ae23
fec7e8e3
fff60793
40e787b3
ffc7f793
00478793
00f70733
00f585b3
01176863
00008067
00050713
ff157ce3
0005c783
00170713
00158593
fef70fa3
ff1768e3
00008067
0045a683
01c5a783
0005af83
0085af03
00c5ae83
0105ae03
0145a303
0185a803
00d72223
0205a683
01f72023
01e72423
01d72623
01c72823
00672a23
01072c23
00f72e23
02470713
40e607b3
fed72e23
02458593
faf2c6e3
f49ff06f
0005c683
00170713
00377793
fed70fa3
00158593
f0078ee3
0005c683
00170713
00377793
fed70fa3
00158593
fc079ae3
f01ff06f
02a5f663
00c587b3
02f57263
00c50733
0e060a63
fff7c683
fff78793
fff70713
00d70023
fef598e3
00008067
00f00793
02c7e863
00050793
fff60693
0c060c63
00168693
00d786b3
0005c703
00178793
00158593
fee78fa3
fed798e3
00008067
00b567b3
0037f793
0a079063
ff060893
ff08f893
01088893
01150833
00058713
00050793
00072683
01070713
01078793
fed7a823
ff472683
fed7aa23
ff872683
fed7ac23
ffc72683
fed7ae23
fcf81ce3
00c67713
011585b3
00f67813
04070e63
00058713
00078893
00300e13
00072303
00470713
40e806b3
0068a023
00d586b3
00488893
fede64e3
ffc80713
ffc77713
00470713
00367613
00e787b3
00e585b3
f39ff06f
00008067
fff60693
00050793
f31ff06f
00008067
00080613
f1dff06f
04c52783
ff010113
00812423
00912223
00112623
01212023
00050413
00058493
02078e63
00249713
00e787b3
0007a503
04050663
00052703
00e7a023
00052823
00052623
00c12083
00812403
00412483
00012903
01010113
00008067
02100613
00400593
0a80a0ef
04a42623
00050793
fa051ae3
00000513
fcdff06f
00100913
00991933
00590613
00261613
00100593
00040513
0780a0ef
fc050ee3
00952223
01252423
f99ff06f
02058063
0045a703
04c52783
00271713
00e787b3
0007a703
00e5a023
00b7a023
00008067
fd010113
03212023
0105a903
01812423
00010c37
02812423
02912223
01312e23
01412c23
01512a23
01612823
02112623
01712623
00058993
00050a13
00060a93
00068413
01458493
00000b13
fffc0c13
0004ab83
000a8593
00448493
018bf533
919f40ef
00850433
000a8593
010bd513
909f40ef
01045793
00f50533
01847433
01051793
008787b3
fef4ae23
001b0b13
01055413
fb2b4ee3
02040263
0089a783
04f95863
00490793
00279793
00f987b3
0087a223
00190913
0129a823
02c12083
02812403
02412483
02012903
01812a03
01412a83
01012b03
00c12b83
00812c03
00098513
01c12983
03010113
00008067
0049a583
000a0513
00158593
e39ff0ef
00050493
04050c63
0109a603
00c98593
00c50513
00260613
00261613
bd1ff0ef
0049a703
04ca2783
00271713
00e787b3
0007a703
00e9a023
0137a023
00490793
00048993
00279793
00f987b3
0087a223
00190913
0129a823
f65ff06f
000256b7
00025537
ef868693
00000613
0b500593
f7850513
64d090ef
fe010113
00812c23
01212823
00058413
00050913
00900593
00868513
00912a23
01312623
01412423
00112e23
01512223
00068493
00060993
00070a13
fe8f40ef
00900793
0c97d863
00100793
00000593
00179793
00158593
fea7cce3
00090513
d5dff0ef
00050593
0a050a63
00100793
00f52823
01452a23
00900793
0937d663
00940a93
01340a33
000a8413
00044683
00a00613
00090513
fd068693
dedff0ef
00140413
00050593
ff4412e3
ff898413
008a8433
0299d663
413484b3
009404b3
00044683
00a00613
00090513
fd068693
db9ff0ef
00140413
00050593
fe8492e3
01c12083
01812403
01412483
01012903
00c12983
00812a03
00412a83
00058513
02010113
00008067
00a40413
00900993
fa5ff06f
00000593
f45ff06f
000256b7
00025537
ef868693
00000613
0ce00593
f7850513
515090ef
ffff0737
00e57733
00050793
00000513
00071663
01079793
01000513
ff000737
00e7f733
00071663
00850513
00879793
f0000737
00e7f733
00071663
00450513
00479793
c0000737
00e7f733
00071663
00250513
00279793
0007ca63
40000737
00e7f7b3
00150513
00078463
00008067
02000513
00008067
00052783
00050713
0077f693
02068463
0017f693
00000513
04069e63
0027f693
0a068863
0017d793
00f72023
00100513
00008067
01079693
0106d693
00000513
06068e63
0ff7f693
06068063
00f7f693
04068263
0037f693
02068463
0017f693
00069c63
0017d793
00150513
00079663
02000513
00008067
00f72023
00008067
0027d793
0017f693
00250513
fe0696e3
fd5ff06f
0047d793
0037f693
00450513
fa069ee3
fddff06f
0087d793
00f7f693
00850513
fa0690e3
fddff06f
0107d793
0ff7f693
01000513
f80692e3
fddff06f
0027d793
00f72023
00200513
00008067
04c52783
ff010113
00812423
00912223
00112623
00050413
00058493
02078c63
0047a503
06050263
00052703
00e7a223
00c12083
00812403
00100793
00952a23
00052623
00f52823
00412483
01010113
00008067
02100613
00400593
3dd090ef
04a42623
00050793
fa051ce3
000256b7
00025537
ef868693
00000613
14000593
f7850513
335090ef
01c00613
00100593
00040513
3a5090ef
fc050ae3
00100793
00f52223
00200793
00f52423
f85ff06f
fb010113
03312e23
03812423
01062983
0105ac03
04812423
03412c23
04112623
04912223
05212023
03512a23
03612823
03712623
03912223
03a12023
01b12e23
00058a13
00060413
013c4c63
00098713
00058413
000c0993
00060a13
00070c13
00842783
00442583
01898bb3
0177a7b3
00f585b3
a09ff0ef
00a12623
20050a63
00c12783
002b9a93
01478b13
015b0ab3
000b0793
015b7863
0007a023
00478793
ff57ece3
014a0a13
002c1c13
01440793
018a0733
00299993
00f12423
00e12023
013789b3
14ea7863
00400713
01540793
00e12223
1af9f263
000104b7
fff48493
01c0006f
0107dc13
0a0c1063
00012783
004a0a13
004b0b13
10fa7e63
000a2783
0097fd33
fe0d00e3
00812c03
000b0c93
00000413
000c2d83
000ca903
000d0593
009df533
b9cf40ef
009977b3
00f507b3
000d0593
010dd513
00878433
01095913
b80f40ef
01045793
01250533
00f50533
00947433
01051793
0087e7b3
004c0c13
00fca023
004c8c93
01055413
fb3c64e3
00412783
00fb07b3
0087a023
000a2783
0107dc13
f60c04e3
000b2403
00812d83
000b0d13
00040913
00000c93
000da503
000c0593
01095913
00957533
b14f40ef
012507b3
01978cb3
00947433
010c9613
00866633
00cd2023
002dd503
004d2903
000c0593
aecf40ef
00997633
010cd793
00c50433
00f40433
004d8d93
004d0d13
01045c93
fb3de4e3
00412783
004a0a13
00fb07b3
0087a023
00012783
004b0b13
eefa66e3
01704863
0180006f
fffb8b93
000b8863
ffcaa783
ffca8a93
fe0788e3
00c12783
04c12083
04812403
0177a823
04412483
04012903
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
00078513
05010113
00008067
408987b3
feb78793
ffc7f793
00478793
00f12223
e4dff06f
000256b7
00025537
ef868693
00000613
15d00593
f7850513
061090ef
fe010113
00812c23
01212823
01312623
00112e23
00912a23
00367793
00060413
00050993
00058913
0a079e63
40245413
06040663
0489a483
0c048a63
00147793
02079063
40145413
04040a63
0004a503
06050663
00050493
00147793
fe0784e3
00048613
00090593
00098513
ce9ff0ef
06090663
00492703
04c9a783
40145413
00271713
00e787b3
0007a703
00e92023
0127a023
00050913
fa041ae3
01c12083
01812403
01412483
00c12983
00090513
01012903
02010113
00008067
00048613
00048593
00098513
c8dff0ef
00a4a023
00052023
00050493
f81ff06f
00050913
f65ff06f
fff78793
00024737
f5870713
00279793
00f707b3
0007a603
00000693
f9cff0ef
00050913
f25ff06f
00100593
00098513
ebcff0ef
00050493
02050063
27100793
00f52a23
00100793
00f52823
04a9a423
00052023
f05ff06f
000256b7
00025537
ef868693
00000613
14000593
f7850513
708090ef
fe010113
01412423
0105aa03
0085a783
01312623
40565993
01498a33
00812c23
00912a23
01212823
01512223
00112e23
001a0913
00058493
00060413
0045a583
00050a93
0127d863
00179793
00158593
ff27cce3
000a8513
e20ff0ef
10050c63
01450813
03305463
00598993
00299993
01350733
00080793
00478793
fe07ae23
fee79ce3
fec98993
01380833
0104a883
01448793
01f47613
00289893
011788b3
0a060463
02000593
40c585b3
00080313
00000693
0007a703
00430313
00478793
00c71733
00d76733
fee32e23
ffc7a683
00b6d6b3
ff17e0e3
01548793
00400713
00f8ea63
409887b3
feb78793
ffc7f793
00478713
00e80833
00d82023
00068463
00090a13
0044a703
04caa783
01c12083
00271713
00e787b3
0007a703
01452823
01812403
00e4a023
0097a023
01012903
01412483
00c12983
00812a03
00412a83
02010113
00008067
0007a703
00478793
00480813
fee82e23
fb17f6e3
0007a703
00478793
00480813
fee82e23
fd17eee3
f95ff06f
000256b7
00025537
ef868693
00000613
1d900593
f7850513
578090ef
01052703
0105a783
00050813
40f70533
04f71263
00279793
01480813
01458593
00f80733
00f587b3
0080006f
02e87463
ffc72683
ffc7a603
ffc70713
ffc78793
fec686e3
00c6b6b3
40d006b3
0016e513
00008067
00008067
0105a703
01062783
ff010113
00812423
00912223
01212023
00112623
00058493
00060413
40f70933
1af71463
00279693
01458593
01460713
00d587b3
00d70733
0080006f
18f5fc63
ffc7a603
ffc72683
ffc78793
ffc70713
fed606e3
16d66063
0044a583
c2cff0ef
1a050263
0104ae03
01042583
01448493
002e1e93
01440813
00259593
01450613
000108b7
01252623
01d48eb3
00b805b3
00060f13
00048313
00000f93
fff88893
00032783
00082683
004f0f13
0117f733
01f70733
0116ffb3
41f70733
0106d693
0107d793
40d787b3
41075693
00d787b3
01079693
01177733
00e6e733
00480813
feef2e23
00430313
4107df93
fab86ae3
408586b3
feb68693
01540413
0026d693
00000793
0085e463
00269793
00f607b3
00400813
0085e663
00168693
00269813
010484b3
010608b3
05d4fe63
00010837
00088593
00048613
fff80813
00062783
00458593
00460613
0107f6b3
01f686b3
4106d713
0107d793
00e787b3
01079713
0106f6b3
00d76733
fee5ae23
4107df93
fdd666e3
fffe8e93
409e8eb3
ffcefe93
01d887b3
00071a63
ffc7a703
fffe0e13
ffc78793
fe070ae3
00c12083
00812403
01c52823
00412483
00012903
01010113
00008067
00048793
00100913
00040493
00078413
e95ff06f
fe0946e3
00000913
e89ff06f
00000593
ab0ff0ef
04050263
00c12083
00812403
00100793
00f52823
00052a23
00412483
00012903
01010113
00008067
000256b7
00025537
ef868693
00000613
24000593
f7850513
2f8090ef
000256b7
00025537
ef868693
00000613
23200593
f7850513
2dc090ef
7ff007b7
00b7f5b3
fcc007b7
00f585b3
00000793
00b05663
00078513
00008067
40b005b3
4145d593
01300793
00b7cc63
000807b7
40b7d5b3
00000793
00078513
00008067
fec58593
01e00713
00100793
00b74663
800007b7
00b7d7b3
00000593
00078513
00008067
fe010113
00912a23
01052483
00812c23
01450413
00249493
009404b3
01212823
ffc4a903
01312623
01412423
00090513
00058993
00112e23
d28ff0ef
02000713
40a707b3
00f9a023
00a00793
ffc48a13
08a7d063
ff550513
05447063
ff84a783
04050063
40a706b3
00d7d733
00a91933
00e96933
ff848613
3ff00737
00e96733
00a797b3
02c47263
ff44a603
00d656b3
00d7e7b3
0140006f
00000793
06051463
3ff00737
00e96733
01c12083
01812403
01412483
01012903
00c12983
00812a03
00078513
00070593
02010113
00008067
00b00693
40a686b3
3ff007b7
00d95733
00f76733
00000793
01447663
ff84a783
00d7d7b3
01550513
00a91933
00f967b3
fa9ff06f
00a91933
3ff00737
00e96733
00000793
f95ff06f
fd010113
01512a23
00058a93
00100593
02912223
01312e23
01412c23
02112623
02812423
03212023
00060493
00068a13
00070993
898ff0ef
10050463
00100737
0144d913
fff70793
7ff97913
00050413
0097f7b3
00090463
00e7e7b3
00f12623
060a9263
00c10513
c58ff0ef
00c12703
00100493
00942823
00e42a23
02050793
08090863
bcd90913
00f90933
03500493
012a2023
40f48533
00a9a023
02c12083
00040513
02812403
02412483
02012903
01c12983
01812a03
01412a83
03010113
00008067
00810513
01512423
bf4ff0ef
00c12703
00050793
04050e63
00812603
02000693
40a686b3
00d716b3
00c6e6b3
00a75733
00d42a23
00e12623
00e034b3
00148493
00e42c23
00942823
f6091ce3
00249713
00e40733
01072503
bce78793
00fa2023
b24ff0ef
00549493
40a48533
f69ff06f
00812683
00d42a23
fc1ff06f
000256b7
00025537
ef868693
00000613
30a00593
f7850513
000090ef
fd010113
03212023
00058913
00810593
02112623
02812423
02912223
01312e23
00050993
d69ff0ef
00050493
00058413
00090513
00c10593
d55ff0ef
01092703
0109a783
00c12683
40e787b3
00812703
00579793
40d70733
00e787b3
00050713
02f05e63
01479793
00878433
00058693
00048513
00040593
00070613
6a00f0ef
02c12083
02812403
02412483
02012903
01c12983
03010113
00008067
01479793
40f585b3
fc9ff06f
ff010113
01212023
00112623
00812423
00912223
01700793
00050913
04a7da63
00025737
0d872783
0dc72583
00025737
0e072403
0e472483
00078513
00040613
00048693
064100ef
fff90913
00050793
fe0914e3
00c12083
00812403
00412483
00012903
00078513
01010113
00008067
00024737
00351913
f5870713
01270733
01072783
00c12083
00812403
01472583
00412483
00012903
00078513
01010113
00008067
01062683
fff58593
4055d593
00158593
01460793
00269693
00259593
00d786b3
00b505b3
02d7f863
00050713
0007a803
00478793
00470713
ff072e23
fed7e8e3
40c687b3
feb78793
ffc7f793
00478793
00f50533
00b57863
00450513
fe052e23
feb56ce3
00008067
01052703
4055d613
01450693
02c75263
00271713
00e687b3
04f6f263
ffc7a703
ffc78793
fe070ae3
00100513
00008067
00261793
00f687b3
fee650e3
01f5f593
fc058ce3
0007a603
00100513
00b65733
00b71733
fce602e3
00008067
00000513
00008067
ff010113
00058713
00812423
00912223
00060593
00050413
042594b7
00068613
00070513
00112623
b404a823
f00f30ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
04001737
00050793
9e472503
00058613
00078593
0040006f
fd010113
03212023
02112623
02812423
02912223
01312e23
01412c23
01512a23
01612823
01712623
01812423
00060913
1c058663
00058413
00050993
dc9f40ef
00b90493
01600713
ffc42783
0e977c63
ff84f493
00048713
0e04cc63
0f24ea63
ffc7fa13
ff840a93
12ea5e63
040006b7
44868c13
008c2583
014a8633
00462683
1ec58063
ffe6f593
00b605b3
0045a583
0015f593
14059663
ffc6f693
00da05b3
0ee5d863
0017f793
02079463
ff842b83
417a8bb3
004ba783
ffc7f793
00d786b3
01468b33
36eb5063
00fa0b33
2ceb5263
00090593
00098513
c98f40ef
00050913
04050c63
ffc42783
ff850713
ffe7f793
00fa87b3
28e78663
ffca0613
02400793
30c7ec63
01300713
22c76063
00050793
00040713
00072683
00d7a023
00472683
00d7a223
00872703
00e7a423
00040593
00098513
f25f30ef
00098513
ccdf40ef
01c0006f
01000493
01000713
f124fae3
00c00793
00f9a023
00000913
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00090513
02012903
03010113
00008067
00c62783
00862703
00058a13
00f72623
00e7a423
004aa783
409a06b3
00f00613
0017f793
014a8733
06d66c63
00fa67b3
00faa223
00472783
0017e793
00f72223
00098513
c35f40ef
00040913
f81ff06f
0017f793
ee0796e3
ff842b83
417a8bb3
004ba783
ffc7f793
ed1ff06f
02812403
02c12083
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00060593
03010113
b44f406f
0097e7b3
00faa223
009a85b3
0016e693
00d5a223
00472783
00858593
00098513
0017e793
00f72223
e01f30ef
f75ff06f
ffc6f693
00da0633
01048593
0eb65063
0017f793
e4079ee3
ff842b83
417a8bb3
004ba783
ffc7f793
00d786b3
01468b33
e2bb4ce3
00cba783
008ba703
ffca0613
02400693
00f72623
00e7a423
008b8913
26c6e063
01300713
00090793
02c77263
00042703
01b00793
00eba423
00442703
00eba623
24c7e663
00840413
010b8793
00042703
00e7a023
00442703
00e7a223
00842703
00e7a423
009b8733
409b07b3
00ec2423
0017e793
00f72223
004ba783
00098513
0017f793
0097e7b3
00fba223
ae9f40ef
e39ff06f
00042683
01b00713
00d52023
00442683
00d52223
18c76663
00840713
00850793
dcdff06f
009a8ab3
409607b3
015c2423
0017e793
00faa223
ffc42783
00098513
00040913
0017f793
0097e7b3
fef42e23
a91f40ef
de1ff06f
ffc52783
ffc7f793
00fa0a33
e19ff06f
00cba783
008ba703
ffca0613
02400693
00f72623
00e7a423
008b8913
10c6e063
01300713
00090793
02c77c63
00042703
01b00793
00eba423
00442703
00eba623
10c7fc63
00842783
00fba823
00c42783
00fbaa23
0ad60663
01040413
018b8793
00042703
000b0a13
000b8a93
00e7a023
00442703
00e7a223
00842703
00090413
00e7a423
d91ff06f
00040593
f98fe0ef
d0dff06f
00c62783
00862703
02400693
ffca0613
00f72623
00e7a423
008ba703
00cba783
008b8913
00f72623
00e7a423
04c6ee63
01300713
00090793
f8c77ae3
00042703
01b00793
00eba423
00442703
00eba623
06c7fa63
00842703
02400793
00eba823
00c42703
00ebaa23
f4f61ee3
01042703
020b8793
01840413
00ebac23
ffc42703
00ebae23
f49ff06f
00040593
00090513
f00fe0ef
00090413
000b0a13
000b8a93
ce1ff06f
00842703
00e52423
00c42703
00e52623
00f60e63
01040713
01050793
c31ff06f
00840413
010b8793
f01ff06f
01042683
01840713
01850793
00d52823
01442683
00d52a23
c09ff06f
00040593
00090513
e9cfe0ef
dddff06f
00842783
00fba823
00c42783
00fbaa23
00d60863
01040413
018b8793
da5ff06f
01042703
020b8793
01840413
00ebac23
ffc42703
00ebae23
d89ff06f
fe010113
01212823
0005a903
00812c23
00912a23
00112e23
01312623
01412423
00058413
00050493
04090263
00092983
02098863
0009aa03
000a0e63
000a2583
00058463
fbdff0ef
000a0593
00048513
aadf30ef
00098593
00048513
aa1f30ef
00090593
00048513
a95f30ef
00040593
01812403
01c12083
01012903
00c12983
00812a03
00048513
01412483
02010113
a6df306f
040017b7
9e47a783
10a78a63
04c52583
fe010113
00912a23
00112e23
00812c23
01212823
01312623
00050493
04058063
00000913
08000993
012587b3
0007a403
00040e63
00040593
00042403
00048513
a19f30ef
fe0418e3
04c4a583
00490913
fd391ce3
00048513
a01f30ef
0404a583
00058663
00048513
9f1f30ef
1484a403
02040063
14c48913
01240c63
00040593
00042403
00048513
9d1f30ef
fe8918e3
0544a583
00058663
00048513
9bdf30ef
0384a783
04078663
03c4a783
00048513
000780e7
2e04a403
02040c63
00042583
00058663
00048513
e95ff0ef
00040593
01812403
01c12083
01012903
00c12983
00048513
01412483
02010113
96df306f
01c12083
01812403
01412483
01012903
00c12983
02010113
00008067
00008067
0005c803
05e00793
00050613
06f80863
00158513
00000693
00000593
00060793
10060713
00d78023
00178793
fee79ce3
04080263
0015c713
02d00313
05d00893
010607b3
00e78023
00054783
00150693
04678063
01178c63
00078863
00078813
00068513
fddff06f
00008067
00068513
00008067
fff50513
00008067
0015c803
00258513
00100693
00100593
f91ff06f
00154583
05158263
0505c063
00250513
00080793
00178793
00f606b3
00e68023
feb7cae3
00180693
00000793
00b84663
00f68833
f85ff06f
410585b3
fff58793
00f68833
f75ff06f
02d00813
00068513
f61ff06f
000257b7
0e87a503
00008067
ff010113
00912223
800004b7
00812423
00112623
fff4c493
00060413
00062023
00b4f6b3
7ff00637
00058793
00050713
06c6d063
00a6e8b3
04088c63
00c5f633
00058813
00000893
02061263
000257b7
0f47a683
0f07a603
65c0f0ef
00050713
00058813
00b4f6b3
fca00893
4146d693
801007b7
fff78793
c0268693
00f87833
011686b3
3fe007b7
00f867b3
00d42023
00c12083
00812403
00412483
00070513
00078593
01010113
00008067
f6010113
08c10e93
08f12a23
80000337
ffff07b7
00058e13
fff34313
08d12623
20878793
00810593
000e8693
06112e23
00f12a23
08e12823
09012c23
09112e23
01c12423
01c12c23
00612e23
00612823
01d12223
5bc040ef
00812783
00078023
07c12083
0a010113
00008067
00050e13
04001537
f6010113
9e452503
08810e93
08f12a23
80000337
ffff07b7
fff34313
08c12423
08d12623
20878793
00058613
000e8693
00810593
06112e23
00f12a23
08e12823
09012c23
09112e23
01c12423
01c12c23
00612e23
00612823
01d12223
540040ef
00812783
00078023
07c12083
0a010113
00008067
00b567b3
0037f793
08079263
0005a703
7f7f86b7
f7f68693
00d777b3
00d787b3
00e7e7b3
00d7e7b3
fff00613
06c79e63
00050613
fff00813
00e62023
0045a703
00458593
00460613
00d777b3
00d787b3
00e7e7b3
00d7e7b3
ff0780e3
0005c783
0015c703
0025c683
00f60023
00078a63
00e600a3
00070663
00d60123
00069463
00008067
000601a3
00008067
00050793
0005c703
00178793
00158593
fee78fa3
fe0718e3
00008067
00050613
fb1ff06f
00b567b3
0037f793
00050713
06079863
00300793
06c7f463
feff0337
808088b7
eff30313
08088893
00300e13
0005a683
006687b3
fff6c813
0107f7b3
0117f7b3
02079e63
00d72023
ffc60613
00470713
00458593
fcce6ce3
00158593
00170793
02060463
fff5c683
fff60813
fed78fa3
00068e63
00078713
00080613
00158593
00170793
fe0610e3
00008067
00c70733
00080a63
00178793
fe078fa3
fee79ce3
00008067
00008067
f4010113
000257b7
0b312623
9207a983
0a812c23
00050413
00098513
0a912a23
0b212823
0b412423
0b512223
09912a23
00060a13
00058c93
00068a93
0a112e23
0b612023
09712e23
09812c23
09a12823
09b12623
06012823
b35f40ef
000247b7
00050613
00000913
00000493
000c8713
02d00513
08078693
06e12623
00074783
00070b93
00f56a63
00279593
00d585b3
0005a583
00058067
00012223
03000713
00000d93
1ce78a63
02f00713
00078493
44f77e63
000b8513
00000d13
00000c13
00000b13
03900713
00800813
02f00593
10974c63
0f684e63
002c1693
01868c33
001c1c13
00fc0c33
fd0c0c13
00150513
06a12623
00054483
001b0b13
00048793
fc95c8e3
00098593
00c12423
314090ef
00812603
000b0793
40051e63
06c12703
00000a93
00c70733
06e12623
00074483
fd048613
00900713
3cc76663
06c12303
00150513
00060493
640610e3
00130713
06e12623
00134483
fd9ff06f
00100793
00f12223
00170b93
07712623
00174783
f20796e3
000a0463
019a2023
00000a93
00000993
0bc12083
0b812403
0b412483
0b012903
0a812a03
0a012b03
09c12b83
09812c03
09412c83
09012d03
08c12d83
000a8513
00098593
0a412a83
0ac12983
0c010113
00008067
00170713
eadff06f
002d1693
01a68d33
001d1d13
00fd0d33
fd0d0d13
f09ff06f
00098593
00c12423
230090ef
0a051c63
06c12783
00812603
00c787b3
06f12623
0007c483
000b0463
7490006f
03000713
64e494e3
00100713
40f70733
03000693
00e78533
00178793
06f12623
0007c483
fed488e3
fcf48793
00800713
2af76a63
06c12b83
fd048493
00150a93
000b8313
00100b13
00000793
002c1713
01870733
00171713
00e48c33
00000513
ed9ff06f
001bc783
05800693
001b8b13
0df7f793
4ad784e3
07612623
000b4783
000b0b93
001b0b13
fee788e3
2a078463
00100d93
e01ff06f
000b0793
00000513
00000a93
00000613
fdf4f713
04500693
00000993
08d71263
00ab6733
01b76733
ea0700e3
06c12c83
02b00713
001c8693
06d12623
001cc483
40e488e3
02d00713
00000593
00e49a63
00100593
002c8713
06e12623
002cc483
fd048713
00900693
78e6e463
03000713
02e49063
06c12703
03000693
00170713
06e12623
00074483
00170713
fed48ae3
fcf48713
00800693
00000993
14e6fae3
080b1a63
00ade533
1e051a63
e0061ee3
06900793
2cf486e3
0697c663
04900793
2cf480e3
04e00793
e0f490e3
000255b7
fd858593
06c10513
51d080ef
de0506e3
06c12703
02800793
00074703
6ef702e3
00025537
e3c50513
06c090ef
00050a93
00058993
000a0663
06c12783
00fa2023
00412783
dc0782e3
800007b7
0137c9b3
db9ff06f
06e00793
faf482e3
da0a10e3
da1ff06f
41598733
00e12623
00079463
000b0793
01000713
000b0c93
01675463
01000c93
000c0513
00f12423
06c100ef
00900713
00812783
00050913
00058493
05675a63
ff7c8713
000246b7
f6868693
00371713
00d70733
00072603
00472683
78d0e0ef
00050913
000d0513
00058493
028100ef
00050613
00058693
00090513
00048593
5590d0ef
00812783
00050913
00058493
00f00713
0f674063
415986b3
1a0682e3
41598633
38c058e3
01600693
48c6dce3
02500693
419b0cb3
41598633
416686b3
00cc8cb3
0cc6c063
41670b33
000249b7
f6898993
003b1793
013787b3
0007a503
0047a583
00090613
00048693
6fd0e0ef
00c12783
416787b3
00379793
013787b3
0007a603
0047a683
6e10e0ef
00050a93
00058993
ebdff06f
00000793
00000a93
00000b13
00100613
db5ff06f
00098593
000b8513
00c12423
709080ef
00812603
3e0504e3
00000793
00000d13
00000c13
00000b13
00000513
00000a93
00000613
00000993
e09ff06f
00000a93
00000993
e61ff06f
419b0cb3
41598733
00ec8cb3
5d905063
00fcf713
02070c63
000246b7
f6868693
00371713
00d70733
00072503
00472583
00090613
00048693
00f12423
6390e0ef
00812783
00050913
00058493
ff0cfc93
760c9c63
02012623
000c0713
000b0693
00078613
000b8593
00040513
e6dfd0ef
02a12823
1a050ae3
00025737
10072683
10472703
00c12583
02d12023
02e12223
00025737
0d872683
0dc72703
fff5c793
04d12823
04e12a23
00025737
12072683
12472703
41f7d793
04d12c23
04e12e23
00025737
11072683
11472703
03412a23
04d12023
04e12223
00025737
11872683
11c72703
02c12a03
413a89b3
04e12623
00f5f7b3
41f5d713
04d12423
00e9fcb3
00f12823
00000c13
00000b13
00050a93
004aa583
00040513
b7dfd0ef
00050b93
20050863
010aa603
00ca8593
00c50513
00260613
00261613
915fd0ef
07810713
07410693
00048613
00090593
00040513
a79fe0ef
06a12823
03212423
00912e23
1a050863
00100593
00040513
ffdfd0ef
00050b13
1a050e63
07412783
3807c263
01012703
019789b3
07812583
414787b3
03600d93
00b787b3
fff78793
c0200613
40bd8db3
20c7d263
40f60633
01f00593
40cd8db3
34c5ce63
00100793
00c797b3
00f12a23
00012c23
01b707b3
01b98db3
00fa0d33
00098713
013dd463
000d8713
00ed5463
000d0713
00e05863
40ed8db3
40ed0d33
40e989b3
0b904c63
0fb04e63
00c12783
18f04263
11a04863
01305e63
000b0593
00098613
00040513
c00fe0ef
00050b13
10050663
07012583
000b8613
00040513
dd0fe0ef
00050c13
0e050a63
00c52783
000b0593
00052623
00f12423
d5cfe0ef
300544e3
1c0508e3
000b0593
000c0513
ac1fe0ef
02012603
02412683
00050d13
00058993
3190e0ef
12a04e63
00812783
2a079663
46090863
00100793
00f91463
4e048ae3
3ff006b7
00000713
bff007b7
00012a23
00d12c23
1440006f
000b0593
000c8613
00040513
a08fe0ef
00050b13
06050663
07012603
00050593
00040513
f45fd0ef
04050c63
07012583
00a12423
00040513
a55fd0ef
00812703
06e12823
f1b056e3
07012583
000d8613
00040513
b18fe0ef
06a12823
ee051ae3
03412a03
0240006f
000b8593
000d0613
00040513
af8fe0ef
00050b93
ee0510e3
03412a03
07012503
02200793
00f42023
00000a93
7ff009b7
00050593
00040513
9edfd0ef
000b8593
00040513
9e1fd0ef
000b0593
00040513
9d5fd0ef
03012583
00040513
9c9fd0ef
000c0593
00040513
9bdfd0ef
ad9ff06f
01012603
000b8593
00040513
930fe0ef
00050b93
f8050ae3
e7a056e3
f75ff06f
00100793
00012c23
00f12a23
e15ff06f
000257b7
0fc7a683
0f87a603
000d0513
00098593
2a90e0ef
00812683
00a12a23
00b12c23
00050713
00058793
00069663
800006b7
00b6c7b3
7ff00337
0064fd33
7fe006b7
00070993
00078d93
14dd0863
060a0e63
06a007b7
07a7ea63
000257b7
1087a603
10c7a683
01412703
01812783
00070513
00078593
1610e0ef
04a04263
01412d83
01812783
000d8513
00078593
1b50f0ef
00051463
00100513
2cd0f0ef
00812783
00a12a23
00b12c23
00050993
68079c63
800007b7
00b7c7b3
00078d93
06b007b7
01b787b3
41a78db3
00090513
00048593
dbcfe0ef
00050613
00058693
00098513
000d8593
1d50e0ef
00090613
00048693
7b80d0ef
00058493
00050913
00058993
000a1863
7ff007b7
00f9f7b3
46fd0863
07012583
00040513
869fd0ef
000b8593
00040513
85dfd0ef
000b0593
00040513
851fd0ef
000c0593
00040513
845fd0ef
c15ff06f
01012703
000c8993
40f70733
c7dff06f
be200613
40f607b3
00100d13
00fd17b3
00f12c23
00100793
00f12a23
c9dff06f
3ff006b7
00000713
3ff007b7
00012a23
00d12c23
eadff06f
07912623
00000993
8a9ff06f
fcb006b7
00d484b3
00090513
00048593
02f12e23
02e12c23
cdcfe0ef
03812703
03c12783
00070613
00078693
0f50e0ef
00090613
00048693
6d80d0ef
7ff00337
00b37733
7ca007b7
00050913
20f76c63
01c12783
fff30313
00679863
02812703
fff00793
d6f70ce3
7ff004b7
fff48493
fff00913
f05ff06f
a80c84e3
41900cb3
00fcf713
02070c63
000246b7
f6868693
00371713
00d70733
00072603
00472683
00090513
00048593
00f12423
6410d0ef
00812783
00050913
00058493
404cdc93
a40c80e3
01f00713
0d974463
010cf713
02e12623
00070663
06a00713
02e12623
00024d37
00090813
00048713
178d0d13
00000613
00078d93
001cf793
02078263
000d2603
004d2683
00080513
00070593
0110e0ef
00050813
00058713
00100613
401cdc93
008d0d13
fc0c98e3
000d8793
00060663
00080913
00070493
02c12703
02070863
0144d693
7ff6f693
06b00713
40d70733
00e05e63
01f00613
06e65ae3
03400613
00000913
06e65ce3
037004b7
00090513
00048593
00000613
00000693
00f12423
5480e0ef
00812783
96051ce3
02200793
00f42023
00000a93
00000993
f68ff06f
00c49793
b8079ee3
05012603
05412683
000d0513
00098593
6800e0ef
4e054e63
000257b7
0f87a603
0fc7a683
000d0513
00098593
7480e0ef
800007b7
00050713
00a12a23
00b12c23
00b7c7b3
cadff06f
06c12303
fd048993
02f00713
00130693
06d12623
00134483
03900813
02f00893
1a975e63
02984663
00299713
01370733
00068e13
00168693
00171713
06d12623
00970733
001e4483
fd070993
fc98cce3
406686b3
00800713
18d75263
000059b7
e1f98993
e4058663
413009b3
e44ff06f
035004b7
00b484b3
00048993
cf9ff06f
13400713
25974e63
404cdd13
00100713
65a75063
00024db7
00048713
058d8693
00000c93
00040493
00090813
000c8413
00d12423
058d8d93
00000613
00100313
00f12823
00070593
00070c93
001d7713
02070063
000da603
004da683
00080513
64c0e0ef
00050813
00100613
00100313
401d5d13
00140413
008d8d93
fc6d18e3
000c8693
01012783
00040c93
00048413
00068493
00060663
00080913
00058493
00f12823
00812783
003c9713
00090613
00e78cb3
000ca503
004ca583
fcb00737
00970733
00070693
5e40e0ef
7ff004b7
00b4f733
7ca006b7
00050913
18e6e263
7c9006b7
01012783
46e6f063
fff48493
fff00913
02012623
f98ff06f
00012223
b48ff06f
00090a93
00048993
d88ff06f
000255b7
fcc58593
06c10513
268080ef
b2050c63
06c12783
000255b7
fd058593
fff78793
06c10513
06f12623
248080ef
00051863
06c12783
00178793
06f12623
00000a93
7ff009b7
d3cff06f
00005737
e1f70713
e93750e3
00070993
e79ff06f
01812d03
01412d83
000d0593
000d8513
6580f0ef
72c0f0ef
00050613
00058693
000d8513
000d0593
3e10e0ef
00812703
00c99793
00c7d793
01276733
00f767b3
00050d13
00058993
02079863
05812603
05c12683
4040e0ef
b2055ee3
03412a03
07012503
00090a93
00048993
9a5ff06f
00000593
c00ff06f
04012603
04412683
3d80e0ef
fc054ce3
04812603
04c12683
000d0513
00098593
2dc0e0ef
aea05ce3
fbdff06f
00412783
00024637
000a8813
07010713
07410693
15060613
06c10593
00040513
0e1070ef
00757a93
00050993
de0a8663
00600793
10fa9263
a00a0a63
016a2023
00000a93
00000993
a0cff06f
02200793
00f42023
ee9ff06f
00100693
001b0713
00aa8ab3
54d50e63
01650533
000b0693
00800813
fff50593
01000893
00070b13
02d86263
002c1693
01868c33
001c1c13
02b70463
00170713
000b0693
00070b13
fed872e3
fee8c6e3
002d1693
01a68d33
001d1d13
fddff06f
00050b13
00800713
a6b75863
01000713
00000513
95674863
002d1713
01a70733
00171713
00e60d33
93cff06f
fea00713
415986b3
d2e6cc63
413a87b3
00024737
f6870713
00379793
00e787b3
0007a603
0047a683
00090513
00048593
1510d0ef
00050a93
00058993
b60ff06f
00058793
00078d93
971ff06f
00000513
9d8ff06f
07012603
00060e63
03500593
07810513
b4cfe0ef
07012583
00040513
a0cfd0ef
00500793
07412683
0357ee63
00024737
002a9793
13870713
00e787b3
0007a783
00078067
07c12483
fff00737
43368793
fff70713
07812903
00e4f4b3
01479793
00f4e4b3
0089f993
00090a93
d40988e3
800009b7
0099e9b3
ad0ff06f
800004b7
fff4c493
fff00913
fddff06f
7ff004b7
fd5ff06f
07812903
07c12483
fc9ff06f
06c12783
00000c13
00000d13
00c787b3
06f12623
0007c483
8f4ff06f
00c12783
00024737
f6870713
00379793
00e787b3
0007a503
0047a583
00090613
00048693
2800e0ef
00050a93
00058993
a5cff06f
000b0793
00000a93
fd1fe06f
3fe006b7
00000713
bfe007b7
00012a23
00d12c23
fccff06f
00812683
00100737
fff70713
03412a03
02812a83
01c12983
00e4f7b3
1a068c63
26e78263
01812783
1a078c63
00f4fcb3
060c8c63
00812783
1c078663
00090513
00048593
dddfd0ef
02c12783
00050693
00058713
02078c63
0144d613
7ff67613
06b00793
40c787b3
02f05263
3ff00737
01479793
00e787b3
00078693
00000613
1cc0e0ef
00050693
00058713
00068613
00090513
00048593
00070693
7a10c0ef
00050a93
00058993
02c12783
04078663
000257b7
1287a603
12c7a683
000a8513
00098593
1880e0ef
00a5e7b3
00050a93
00058993
07012503
e4079463
02200793
00f42023
e3cff06f
035004b7
00b484b3
02012623
b3cff06f
07012503
e24ff06f
000245b7
07810613
16458593
06c10513
659070ef
00500793
00f50463
904ff06f
07c12783
7ff009b7
07812a83
00f9e9b3
904ff06f
00812783
03412a03
02812a83
0127e933
01c12983
f60910e3
00c49793
f4079ce3
7ff007b7
00f4f7b3
06b00737
f4f774e3
014c2783
00079863
010c2703
00100793
f2e7dae3
000c0593
00100613
00040513
871fd0ef
000b0593
00050c13
9f5fd0ef
f0a05ae3
02c12783
12078e63
7ff007b7
00f4f7b3
06b00737
12f74663
03700737
eef74ee3
07012483
02200793
00f42023
00048513
00000a93
00000993
d50ff06f
0127e7b3
e40796e3
fbdff06f
01412783
0127fd33
ec0d00e3
e49ff06f
00024737
05870713
00000c93
00e12423
a41ff06f
00090513
00048593
c15fd0ef
02c12783
00050693
00058713
10078463
0144d613
7ff67613
06b00793
40c787b3
02f05263
3ff00737
01479793
00e787b3
00078693
00000613
0040e0ef
00050693
00058713
00068613
00090513
00070693
00048593
6b40e0ef
00000613
00000693
00050a93
00058993
5810d0ef
e2051ae3
f39ff06f
02c12783
fff00713
02078263
7ff007b7
00f4f7b3
06a006b7
00f6ea63
0147d793
06b00693
40f687b3
00f71733
d6e91ae3
7ff007b7
fff78793
0af48663
7ff009b7
0134f9b3
001007b7
00000a93
00f989b3
dd5ff06f
7ff009b7
fff007b7
0134f9b3
00f989b3
001007b7
fff78793
fff00a93
00f9e9b3
db1ff06f
fff00693
00e69733
01277933
f94ff06f
04b00713
40d706b3
fff00713
00d71733
009774b3
f7cff06f
00068613
00048593
00070693
00090513
5e40e0ef
00000613
07012483
00000693
00050a93
00058993
4ad0d0ef
00050793
00048513
bc079463
e61ff06f
03412a03
e55ff06f
fff00793
f4f91ae3
b9cff06f
000b0593
00070b13
af5ff06f
040016b7
85068693
afdfe06f
04001737
00050793
9e472503
00060693
00058613
00078593
ae1fe06f
04001737
00050793
9e472503
040016b7
00058613
85068693
00078593
ac1fe06f
fd010113
01412c23
04001a37
00050793
9e4a2503
00060693
00058613
00078593
02812423
02912223
02112623
03212023
01312e23
01512a23
01612823
01712623
a7dfe0ef
00050613
00058693
00050493
00058413
4ed0e0ef
0c051263
00040593
00048513
398120ef
000257b7
1387ab03
800009b7
fff9c993
01357ab3
00050913
000b0593
000a8513
138120ef
06051063
000b0593
000a8513
070120ef
04a05863
000257b7
1307ab03
1347ab83
01347433
00048513
00040593
000b0613
000b8693
4810e0ef
00051e63
00048513
00040593
000b0613
000b8693
4c90d0ef
00a04863
9e4a2783
02200713
00e7a023
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00c12b83
00090513
02012903
03010113
00008067
00025537
e3c50513
00045a63
e9cfe0ef
80000937
00a94933
fb9ff06f
02812403
02c12083
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
03010113
e64fe06f
fd010113
01412c23
04001a37
00050793
9e4a2503
040016b7
00058613
85068693
00078593
02812423
02912223
02112623
03212023
01312e23
01512a23
01612823
01712623
915fe0ef
00050613
00058693
00050493
00058413
3850e0ef
0c051263
00040593
00048513
230120ef
000257b7
1387ab03
800009b7
fff9c993
01357ab3
00050913
000b0593
000a8513
7d1110ef
06051063
000b0593
000a8513
709110ef
04a05863
000257b7
1307ab03
1347ab83
01347433
00048513
00040593
000b0613
000b8693
3190e0ef
00051e63
00048513
00040593
000b0613
000b8693
3610d0ef
00a04863
9e4a2783
02200713
00e7a023
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00c12b83
00090513
02012903
03010113
00008067
00025537
e3c50513
00045a63
d34fe0ef
80000937
00a94933
fb9ff06f
02812403
02c12083
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
03010113
cfcfe06f
fe010113
00058813
040017b7
00812c23
00060593
00050413
00068613
85078793
00010713
00000693
00080513
00112e23
7ac000ef
00012783
01c12083
00040513
00f42023
00412783
00f42223
00812783
00f42423
00c12783
00f42623
01812403
02010113
00008067
fe010113
040017b7
00812c23
00050413
9e47a503
00010713
00068793
00000693
00112e23
750000ef
00012783
01c12083
00040513
00f42023
00412783
00f42223
00812783
00f42423
00c12783
00f42623
01812403
02010113
00008067
fe010113
040017b7
00812c23
00050413
9e47a503
040017b7
85078793
00010713
00000693
00112e23
6f0000ef
00012783
01c12083
00040513
00f42023
00412783
00f42223
00812783
00f42423
00c12783
00f42623
01812403
02010113
00008067
fa010113
03912a23
00068c93
000246b7
05212823
04112e23
04812c23
04912a23
05312623
05412423
05512223
05612023
03712e23
03812c23
03a12823
03b12623
00b12a23
00a12e23
00c12423
00058913
c0168693
00094483
00090613
00190913
009687b3
0007c783
0087f793
fe0794e3
02d00793
1ef48063
02b00793
0ef48863
fff00793
80000ab7
00f12823
fffaca93
00012c23
0e0c8c63
01000793
1cfc8a63
000c8d93
41fcd993
01012403
000d8613
00098693
00040513
000a8593
2f80c0ef
00050b93
000d8613
00098693
00040513
000a8593
01712623
51d0b0ef
00050c13
00058a13
00000793
00000513
00000593
00900b93
01900b13
fff00d13
fd048413
008bfe63
fbf48693
fc948413
00db7863
f9f48693
0adb6263
fa948413
09945e63
03a78c63
04ba6063
01459463
02ac6c63
06ac0a63
000d8613
00098693
3a0120ef
41f45793
00a40533
00b785b3
00853433
00b405b3
00100793
00190913
fff94483
f9dff06f
fff00793
ff1ff06f
fff00793
80000ab7
00f12823
00012c23
00094483
fffaca93
00260913
f00c98e3
03000793
10f48e63
00a00d93
00000993
00a00c93
f09ff06f
f8ba18e3
00c12703
fff00793
fa8744e3
f81ff06f
fff00713
06e78863
01812703
00070a63
00a03733
40b005b3
40e585b3
40a00533
00812703
00070a63
0e079663
00812783
01412703
00e7a023
05c12083
05812403
05412483
05012903
04c12983
04812a03
04412a83
04012b03
03c12b83
03812c03
03412c83
03012d03
02c12d83
06010113
00008067
01c12703
02200793
00f72023
00812783
08078e63
fff90793
01012503
00f12a23
000a8593
f95ff06f
00100793
00094483
00012823
00260913
80000ab7
00f12c23
e29ff06f
03000793
00f49a63
00094783
05800693
0df7f793
00d78863
01000d93
00000993
e19ff06f
00194483
01000d93
00290913
00000993
01000c93
e01ff06f
00094783
05800713
0df7f793
fce78ee3
00800d93
00000993
00800c93
de1ff06f
00a12823
00058a93
f6dff06f
01012503
000a8593
f11ff06f
d1dff06f
04001737
00050793
9e472503
00060693
00058613
00078593
d01ff06f
04001737
00050793
9e472503
00060693
00058613
00078593
ce5ff06f
fb010113
04112623
04812423
04912223
05212023
03312e23
03412c23
03512a23
03612823
03712623
03812423
03912223
03a12023
01b12e23
00100793
00a12423
10f68a63
02400793
00068c93
00068a13
10d7e263
00024737
00058913
00060993
00058413
c0170713
00044483
00040693
00140413
009707b3
0007c783
0087f793
fe0794e3
02d00793
1af48063
02b00793
10f48863
80000b37
fffb4b13
00012623
100c8c63
01000793
1afc8263
000a0593
000b0513
f99f00ef
00050b93
000a0593
000b0513
f41f00ef
00900d93
fd048793
00050d13
00000713
00000513
01900a93
fff00c13
02fdee63
00078493
0594d263
03870063
fff00713
00ad6c63
10ad0063
000a0593
ed5f00ef
00a48533
00100713
00044483
00140413
fd048793
fcfdf6e3
fbf48793
0cfae463
fc948493
fd94c2e3
fff00793
0cf70863
00c12783
00078463
40a00533
02098063
12071263
0129a023
0140006f
6d8060ef
01600793
00f52023
00000513
04c12083
04812403
04412483
04012903
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
05010113
00008067
80000b37
00012623
00044483
fffb4b13
00268413
ee0c98e3
03000793
08f49263
00044783
05800713
00800a13
0df7f793
00800c93
ece79ce3
00144483
01000a13
00240413
01000c93
ec5ff06f
f9f48793
f4fae0e3
fa948493
ef5ff06f
f09bcae3
f01ff06f
00812703
02200793
000b0513
00f72023
f40988e3
fff40913
000b0513
0129a023
f41ff06f
00100793
00044483
80000b37
00268413
00f12623
e65ff06f
00a00a13
00a00c93
e65ff06f
03000793
01000a13
e4f49ce3
00044783
05800713
0df7f793
e4e794e3
f71ff06f
00050b13
fa9ff06f
d8dff06f
04001737
00050793
9e472503
00060693
00058613
00078593
d71ff06f
04001737
00050793
9e472503
00060693
00058613
00078593
d55ff06f
0076f793
00600713
04f76a63
00024737
00279793
1a070713
00e787b3
0007a783
00078067
000047b7
03e78793
00f60633
01061613
01065613
0045a783
0005a703
00c51423
0107d613
01075593
00e51023
00b51123
00f51223
00c51323
0086f693
00068a63
00855783
ffff8737
00e7e7b3
00f51423
00008067
00051423
00051323
00051223
00051123
00051023
0086f693
fe0682e3
fd1ff06f
7fff87b7
00052023
00052223
00052423
00f52623
0086f693
fc0682e3
fb1ff06f
ffff87b7
fff7c713
00e51423
00f51323
00051023
00051123
00051223
0086f693
f8068ee3
f89ff06f
00000613
f55ff06f
fd010113
02912223
02112623
02812423
00100893
00070493
00078813
07168863
040018b7
9bc88893
0008ae03
0048a303
0088a703
0108a783
00d12c23
01c12623
00612823
00e12a23
00f12e23
00c10693
00410793
00010713
415070ef
00012603
00050413
00050693
00410593
00048513
ea9ff0ef
02c12083
00040513
02812403
02412483
03010113
00008067
040016b7
9bc68693
fbdff06f
fb010113
00024737
03412c23
03a12023
01b12e23
04112623
04812423
04912223
05212023
03312e23
03512a23
03612823
03712623
03812423
03912223
00058a13
00a12623
00c12023
00068d93
00058d13
c0170713
000d4483
000d0693
001d0d13
009707b3
0007c783
0087f793
fe0794e3
02d00793
1cf48263
02b00793
00012423
10f48263
040d8863
01000793
1cfd8063
41fdd993
000d8613
00098693
fff00513
fff00593
6000b0ef
00058713
00050913
000d8613
00098693
fff00513
fff00593
00070b13
3a10b0ef
000d8c93
00a12223
02c0006f
03000793
1af48c63
000257b7
1407a903
1447ab03
00500793
00f12223
00a00c93
00000993
00a00d93
00000793
00000513
00000593
00900a93
01900b93
fff00c13
fd048413
008afe63
fbf48693
fc948413
00dbf863
f9f48693
06dbec63
fa948413
07b45863
03878c63
04bb6063
01659463
02a96c63
05250463
000c8613
00098693
439110ef
41f45793
00a40533
00b785b3
00853433
00b405b3
00100793
001d0d13
fffd4483
f9dff06f
fff00793
ff1ff06f
000d4483
00268d13
ef9ff06f
fb659ee3
00412703
fff00793
fc874ae3
fadff06f
fff00713
06e78663
00812703
00070a63
00a03733
40b005b3
40e585b3
40a00533
00012703
00070863
06079263
00012783
0147a023
04c12083
04812403
04412483
04012903
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
05010113
00008067
00c12703
02200793
fff00513
00f72023
00012783
fff00593
fa0786e3
fffd0a13
f9dff06f
00100793
000d4483
00f12423
00268d13
e3dff06f
03000793
0af49c63
000d4783
05800713
0df7f793
06e79263
00f00793
10000737
001d4483
00f12223
002d0d13
fff00913
fff70b13
01000c93
00000993
01000d93
e71ff06f
000d4783
05800713
0df7f793
fce784e3
00700793
20000737
00f12223
fff00913
fff70b13
00800c93
00000993
00800d93
e3dff06f
01000613
00000693
fff00513
fff00593
3d00b0ef
00058713
00050913
01000613
00000693
fff00513
fff00593
00070b13
1710b0ef
01000c93
00000993
00a12223
df9ff06f
00f00793
10000737
00f12223
fff00913
fff70b13
01000c93
00000993
dd9ff06f
cd9ff06f
04001737
00050793
9e472503
00060693
00058613
00078593
cbdff06f
04001737
00050793
9e472503
00060693
00058613
00078593
ca1ff06f
fb010113
00024737
04812423
05212023
03312e23
03812423
04112623
04912223
03412c23
03512a23
03612823
03712623
03912223
03a12023
01b12e23
00058913
00a12623
00060993
00068c13
00058413
c0170713
00044483
00040693
00140413
009707b3
0007c783
0087f793
fe0794e3
02d00793
14f48e63
02b00793
00000b13
10f48863
020c0a63
01000793
14fc0a63
000c0593
fff00513
fd8f00ef
00050c93
000c0593
fff00513
811f00ef
000c0b93
00050a93
0200006f
03000793
14f48e63
1999acb7
00500a93
999c8c93
00a00b93
00a00c13
00900d13
fd048793
00000713
00000513
01900a13
fff00d93
02fd6e63
00078493
0584d263
03b70063
fff00713
00acec63
0b950463
000b8593
f38f00ef
00a48533
00100713
00044483
00140413
fd048793
fcfd76e3
fbf48793
06fa6863
fc948493
fd84c2e3
fff00793
06f70c63
000b0463
40a00533
00098663
06071e63
0129a023
04c12083
04812403
04412483
04012903
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
05010113
00008067
00044483
00268413
eedff06f
f9f48793
f8fa6ce3
fa948493
f4dff06f
f69ac6e3
f59ff06f
00c12703
02200793
fff00513
00f72023
f80988e3
fff40913
f85ff06f
00044483
00100b13
00268413
ea9ff06f
03000793
08f49263
00044783
05800713
0df7f793
04e79663
10000cb7
00144483
00f00a93
00240413
fffc8c93
01000b93
01000c13
ec1ff06f
00044783
05800713
0df7f793
fce78ae3
20000cb7
00700a93
fffc8c93
00800b93
00800c13
e99ff06f
01000593
fff00513
e28f00ef
00050c93
01000593
fff00513
e60f00ef
01000b93
00050a93
e71ff06f
10000cb7
00f00a93
fffc8c93
01000b93
e5dff06f
d85ff06f
04001737
00050793
9e472503
00060693
00058613
00078593
d69ff06f
04001737
00050793
9e472503
00060693
00058613
00078593
d4dff06f
ff010113
00112623
00812423
00912223
01212023
fff00793
06f58a63
00c65783
03062683
00462703
fdf7f793
00f61623
00060413
0ff5f913
0ff5f493
04068c63
03462783
02f75e63
00042783
fff78713
00e42023
ff278fa3
00442783
00178793
00f42223
00c12083
00812403
00012903
00048513
00412483
01010113
00008067
00060593
4a0040ef
fc0500e3
fff00493
fd5ff06f
01062683
00062783
00068863
00f6f663
fff7c683
04968663
02f42c23
00300793
05240123
02f42a23
04040613
04240693
00100793
00c12083
02e42e23
02c42823
00d42023
00f42223
00812403
00012903
00048513
00412483
01010113
00008067
fff78793
00170713
00f62023
00e62223
f61ff06f
ff010113
00812423
00058413
0305a583
00112623
02058e63
04040793
00f58463
da5f00ef
03c42783
02042823
00f42223
02078063
03842783
00000513
00f42023
00c12083
00812403
01010113
00008067
00c45783
01042703
00042223
0207e793
00e42023
00f41623
fff00513
fd5ff06f
fd010113
01312e23
01912223
00050993
00058c93
00068513
00060593
02812423
01412c23
01512a23
01612823
02112623
02912223
03212023
01712623
01812423
00060a93
00068b13
00070413
bc8f00ef
00050a13
0a050063
00442483
00042583
00050913
04040b93
06a4f263
000c8513
00048613
f14fb0ef
00042783
03042703
00042223
009787b3
00f42023
00090c13
00070593
00098513
009c8cb3
40990933
08070663
01770463
cadf00ef
03c42783
02042823
00f42223
06078a63
03842583
00078493
00b42023
fb27e2e3
00090613
000c8513
eb4fb0ef
00442703
00042783
000b0a13
41270733
012787b3
00e42223
00f42023
02c12083
02812403
02412483
02012903
01c12983
01412a83
01012b03
00c12b83
00812c03
00412c83
000a0513
01812a03
03010113
00008067
00c45783
01042703
009a0533
0207e793
00e42023
00042223
00f41623
000a8593
41850533
af0f00ef
00050a13
f9dff06f
e4010113
1a812c23
1b312623
19912a23
1c010413
1a112e23
1a912a23
1b212823
1b412423
1b512223
1b612023
19712e23
19812c23
19a12823
19b12623
00c59703
e6d42823
00058993
01271693
00050c93
0206c263
0645a683
000025b7
00b76733
ffffe5b7
fff58593
00b6f6b3
00e99623
06d9a223
00064703
00160913
e8e42223
00071463
6c40106f
000246b7
c0168d93
000246b7
1bc68793
000246b7
e6f42623
31468793
000246b7
e6f42423
44c68793
e6042023
e6042e23
00000c13
e6042a23
00000d13
e6042c23
e4f42e23
00ed86b3
0006c683
0086f693
0c069263
02500693
04d71263
00094683
00000a93
00000493
05500613
06800513
06c00593
fdb68793
0ff7f793
00190713
18f66463
e6c42803
00279793
010787b3
0007a783
00078067
00070913
0049a703
12e05a63
0009a703
00074603
fff94683
0ed60c63
e7c42783
00078c63
e7c42783
0007aa03
000a0663
000a0513
fadf00ef
e7842503
e4040113
1bc12083
1b812403
1b412483
1b012903
1ac12983
1a812a03
1a412a83
1a012b03
19c12b83
19812c03
19412c83
19012d03
18c12d83
1c010113
00008067
0049a683
04098493
02d05c63
0009a783
0007c703
00ed8733
00074703
00877713
06070063
0049a683
00178793
00f9a023
fff68693
00d9a223
001d0d13
fcd048e3
0309a583
64058ae3
00958663
000c8513
a0df00ef
03c9a783
0209a823
00f9a223
62078ce3
0389a783
00f9a023
0007c703
00ed8733
00074703
00877713
fa0714e3
00094703
00190913
e8e42223
ea0712e3
f11ff06f
0049a683
00170713
00e9a023
fff68713
00e9a223
00094703
001d0d13
00190913
e8e42223
e6071ce3
ee5ff06f
0309a583
620584e3
04098713
00e58663
000c8513
989f00ef
03c9a703
0209a823
00e9a223
600704e3
0389a703
00e9a023
ea5ff06f
e7c42783
ec0782e3
0007aa03
eb1ff06f
08faf793
e8079ce3
00249793
009784b3
00149493
00d484b3
fd048493
00194683
00070913
e39ff06f
00faf793
fe0788e3
e6dff06f
00faf793
e60792e3
00194683
002aea93
00070913
e15ff06f
e6e42223
200aea93
00011737
b0870793
e6f42023
01000793
e6f42a23
00300913
0049a703
1ee05863
040af713
22070063
00200713
3ee90c63
00300713
00e90ce3
00100713
5ce90a63
00049463
00100493
001af713
010afa13
200700e3
000a0463
1e40106f
e7042783
080afa93
0007a703
00478793
e4f42623
e6e42823
000a9463
2a00106f
f20700e3
08000513
d79f00ef
00050913
52050ae3
e7c42783
e7042683
0067db03
0047d703
00a6a023
72eb7ae3
0007a503
002b1713
00e50533
e7c42703
001b0793
e5242a23
00f71323
e7042783
00f52023
02000793
e4f42c23
04098793
00000b93
00300a93
fff00b13
e4f42823
c99fa0ef
4d7500e3
0009a783
0049a703
fc0b8693
0007c603
008686b3
fff70713
00178793
ecc68c23
00e9a223
00f9a023
001b8b93
015c1863
e9042783
00400713
00e78a63
00800613
00000593
e9040513
c9cf10ef
e9040713
000b8693
e9840613
00090593
000c8513
f91fa0ef
00050c13
45650ae3
600514e3
000a1463
00092023
017d0d33
fff48493
020a1263
e7042783
00078c63
e5442783
e5842703
40f90bb3
402bd793
60e7fee3
00490913
0049a783
00000b93
5cf05ce3
f40494e3
e7042783
00078e63
e5442783
40f905b3
e5842783
4025d713
00f77463
4340106f
e7842783
001a3a13
e6442903
014787b3
e6f42c23
e4c42783
e6f42823
d49ff06f
e6e42223
001aea93
00011737
b0870793
0049a703
e6f42023
00800793
e6f42a23
00300913
e0e04ce3
0309a583
380582e3
04098713
00e58663
000c8513
ee4f00ef
03c9a703
0209a823
00e9a223
360702e3
0389a703
00e9a023
040af713
de0714e3
0009a683
0006c703
00ed8733
00074703
00877713
dc0708e3
04098a13
01c0006f
00d9a023
0006c783
00fd87b3
0007c783
0087f793
da0788e3
0049a783
001d0d13
00168693
fff78793
00f9a223
fcf04ae3
0309a583
2e058ee3
01458663
000c8513
e60f00ef
03c9a783
0209a823
00f9a223
2e0780e3
0389a683
fa9ff06f
00070593
ec040513
cf5fc0ef
e6a42223
040aea93
00100913
d41ff06f
00faf793
b60794e3
00194683
00b69463
7c90006f
001aea93
00070913
b11ff06f
00faf793
b40794e3
00194683
00a69463
7990006f
004aea93
00070913
af1ff06f
e6e42223
00010737
36c70793
e6f42023
e6042a23
00300913
ce5ff06f
e6e42223
001aea93
00200913
cd5ff06f
e6e42223
001aea93
00010737
36c70793
e6f42023
00a00793
e6f42a23
00300913
cb1ff06f
e6e42223
001aea93
040aea93
00000913
c9dff06f
08faf793
ac0792e3
e7c42783
00079463
7b10006f
00194683
080aea93
00070913
a69ff06f
00070913
010af713
b6071ee3
e7042783
008af713
0007a683
00478613
00071463
7990006f
01a68023
e6c42823
b59ff06f
e6e42223
220aea93
c25ff06f
e6e42223
00200913
c31ff06f
e6e42223
00011737
b0870793
e6f42023
00a00793
e6f42a23
00300913
c11ff06f
0154e4b3
a2049ce3
00194683
01000a93
00070913
9e9ff06f
00049463
fff00493
001afa13
010af913
6e0a0263
5e0918e3
e7042783
080afa93
0007aa03
00478b13
6a0a8ae3
b40a06e3
08000513
9a5f00ef
00050b93
160500e3
e7c42783
00aa2023
0067da83
0047d703
38eafee3
0007a503
e7c42783
002a9713
001a8a93
01579323
00e50533
02000793
01452023
e7642823
000b8a93
e4f42c23
0009a703
00074703
00ed8733
00074703
00877713
10071063
04098793
00000b13
e4f42a23
8b9fa0ef
0f6500e3
0009a783
0049a703
fc0b0693
0007c603
008686b3
00178793
fff70713
00f9a023
ecc68c23
00e9a223
00300793
001b0b13
00fc1863
e9042783
00400713
00e78a63
00800613
00000593
e9040513
8b8f10ef
e9040713
000b0693
e9840613
000b8593
000c8513
badfa0ef
fff00793
00050c13
06f506e3
520512e3
000ba023
e5642823
c09f70ef
00050463
0680106f
016d0d33
fff48493
00090463
7b50006f
004b8b93
000a1463
7a90006f
e5842683
415b87b3
4027d713
00000b13
00d76463
1180106f
0049a783
00f04463
7f50006f
0009a783
0007c783
00fd87b3
0007c783
0087f793
00079463
f0049ae3
04091063
000ba023
020a0663
415b85b3
e5842783
4025d713
00170713
00f77c63
000a2503
00458593
ab4fc0ef
00050463
00aa2023
e7842783
00178793
e6f42c23
e6442903
00094703
00190913
e8e42223
fc071863
83dff06f
00049463
fff00493
010af793
001af713
e4f42c23
5c070a63
32079ae3
e7042783
080afa93
0007a703
00478793
e4f42223
e4e42a23
4e0a84e3
94070ae3
08000513
facf00ef
00050a13
76050463
e7c42783
e5442683
0067d903
0047d703
00a6a023
0ee966e3
000106b7
ff668693
74e6e663
e7c42b03
00870713
01071a93
000b2503
010ada93
002a9593
9fcfc0ef
72050663
00ab2023
015b1223
e7c42783
00291713
00190913
01279323
e5442783
00e50533
e5442823
00f52023
02000793
e4f42623
04098793
04001bb7
00000913
00300a93
e4f42423
850b8b93
e98fa0ef
6d250063
0009a783
0049a703
fc090693
0007c603
008686b3
fff70713
00178793
ecc68c23
00e9a223
00f9a023
00190913
015c1863
e8842703
00400793
00f70a63
00800613
00000593
e8840513
e9df00ef
e8840713
00090693
e9840613
000a0593
000c8513
991fa0ef
fff00793
00050c13
00090813
64f50663
7a051a63
000a2023
00000b13
00800613
00000593
e9040513
e7042823
e55f00ef
0e0ba783
000b0613
e9040693
e8040593
000c8513
000780e7
00100793
e7042803
00000b13
00f51463
e8044b03
fc0b0793
00878b33
f00b4783
52078ae3
012d0d33
755c0263
fff48493
e5842783
02079263
e5442783
004a0a13
00078c63
e5042783
e4c42703
40fa0933
40295793
0ae7fee3
0049a783
00000913
72f05663
ee0494e3
e5842783
02079a63
e5442783
000a2023
00078e63
e5042783
40fa05b3
e4c42783
4025d713
00170713
60f76ae3
e7842783
00178793
e6f42c23
e4442783
e6442903
e6f42823
ee0ff06f
fff48713
02600693
00000613
00e6f663
fd948613
02700493
00001837
e7442883
d8080713
e9840b13
fffffbb7
00eaeab3
00000913
000b0a13
47fb8b93
80080813
0009a703
04d00593
00074683
fd568793
0ff7f793
04f5e663
e6842583
00279793
00b787b3
0007a783
00078067
00a00793
0317d863
017afab3
00da0023
001a0a13
0049a783
00170713
fff78793
00f9a223
0ef05e63
00e9a023
fff48493
fa0492e3
e7142a23
100af713
00070663
594b6c63
d56a0663
010af713
12071c63
e6042783
e7442683
00000613
000b0593
000c8513
000a0023
000780e7
e7042783
020af713
00478493
0e071a63
008af713
70071e63
004af713
360700e3
e7042783
0007a703
00a71023
0dc0006f
e5c42783
00189893
017afab3
011788b3
00089883
f5dff06f
600af793
20000593
f6b79ce3
dffafa93
500aea93
01000893
f41ff06f
080af793
f60780e3
f7fafa93
f31ff06f
e5c42783
00189893
011788b3
00089883
00800793
f117cae3
f3dff06f
010af7b3
f00786e3
00089663
200aea93
00800893
400af793
44078063
a7fafa93
ef1ff06f
0309a583
360588e3
04098793
02f58263
000c8513
e4c42c23
e7142a23
f11ef0ef
e5842603
e7442883
000017b7
80078813
03c9a783
0209a823
00f9a223
32078ce3
0389a703
ec5ff06f
e7042783
0007a703
00a72023
e7842783
e6942823
00178793
e6f42c23
416a0a33
012a0a33
014d0d33
e6442903
bb1ff06f
680a1663
e7042783
080afa93
0007aa03
00478b93
3e0a8863
be0a0063
00048513
b8cf00ef
00050913
34050463
e7c42783
00aa2023
0067da83
0047d703
0007a503
02eaea63
000106b7
ff668693
32e6e663
00870713
01071b13
010b5b13
002b1593
de5fb0ef
30050a63
e7c42783
00a7a023
01679223
e7c42783
002a9713
00e50733
001a8a93
01472023
00090593
01579323
00098713
00048693
00100613
000c8513
8c0ff0ef
00050913
440502e3
36957c63
000a2503
00090593
d8dfb0ef
36050463
00aa2023
3600006f
080918e3
e7042783
080afa93
0007aa03
00478793
e6f42823
720a8463
b00a0a63
02000513
ac0f00ef
00050913
26050e63
e7c42b83
00aa2023
006bda83
004bd703
000ba503
34eaf663
e7c42783
002a9713
00e50533
001a8a93
01579323
01452023
02000b93
0009a703
00074683
00dd86b3
0006c683
0086f693
68069863
00090a93
04098813
0049a783
00170693
00d9a023
fff78793
00f9a223
00074783
00190b13
00f90023
000a0663
415b0933
71797063
fff48493
24048c63
0049a783
78f05e63
0009a703
00074783
00fd87b3
0007c783
0087f793
22079c63
000b0913
fa9ff06f
e5842783
56079e63
e7042783
080afa93
0007ab03
00478793
e6f42823
6c0a8e63
a20b0863
02000513
9dcf00ef
00050a13
18050c63
e7c42b83
00ab2023
006bd903
004bd703
000ba503
28e97c63
e7c42783
00291713
00e50533
00190913
01279323
01652023
02000b93
0009a703
00074683
fc068793
008786b3
f006c683
9c068a63
e5842c23
000a0a93
04098913
000b0c13
0380006f
41578b33
00078a13
097b7463
fff48493
0c048063
0049a783
04f05463
0009a703
00074783
fc078793
008787b3
f007c783
0a078063
0049a783
00170693
00d9a023
fff78793
00f9a223
00074703
001a0793
00ea0023
fa0c16e3
00078a13
fb1ff06f
0309a583
02058ae3
01258663
000c8513
c09ef0ef
03c9a783
0209a823
00f9a223
00078ce3
0389a703
00e9a023
f95ff06f
001b9b93
000a8513
000b8593
b6dfb0ef
00050a93
08050863
01650a33
00ac2023
f5dff06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
9d0ff06f
000c0b13
e5842c03
415a04b3
8f5a0063
000a0023
000b0663
00148593
3175e263
e7842783
e6442903
009d0d33
00178793
e6f42c23
998ff06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
e7842783
00078863
00c9d783
0407f793
88078663
e7c42783
0a078ae3
e7c42783
0067d983
0007aa03
02098663
000a0493
00000913
0004a783
00448493
00190913
0007a503
81cf00ef
ffc4a783
0007a023
ff2992e3
fff00793
e6f42c23
850ff06f
c7fafa93
00060663
fff60613
00148493
00190913
aadff06f
415b0ab3
001a8593
015d0d33
000b0913
00090023
fa0a0a63
fb75f863
000a2503
a51fb0ef
fa050263
00aa2023
f9cff06f
00098713
00048693
00100613
000a0593
000c8513
d49fe0ef
00050913
f2050ee3
e7842783
012d0d33
e7742823
00178793
e6442903
e6f42c23
89cff06f
fffa4583
00098613
000c8513
fffa0a13
b99fe0ef
a59ff06f
000106b7
ff668693
f0e6ece3
00870713
01071b13
010b5b13
002b1593
9d1fb0ef
f00500e3
00aba023
016b9223
c8dff06f
000106b7
ff668693
eee6e4e3
00870713
01071a93
010ada93
002a9593
9a1fb0ef
ec0508e3
00aba023
015b9223
d41ff06f
e8842703
00400793
8af71ce3
8b9ff06f
ffe00713
02e51ee3
0049a783
fcf04263
0309a583
54058a63
e4842783
00f58663
000c8513
9c9ef0ef
03c9a783
0209a823
00f9a223
52078a63
0389a783
00f9a023
8a9ff06f
0007a503
f48ff06f
ffe00793
12f51463
0049a783
96f04c63
0309a583
4e058263
e5042783
00f58663
000c8513
97def0ef
03c9a783
0209a823
00f9a223
4c078263
0389a783
00f9a023
9fcff06f
e5442503
00371593
8e5fb0ef
e4a42a23
e00504e3
e5842783
e7042703
01750933
00179793
00a72023
e4f42c23
9bcff06f
000106b7
ff668693
dee6e4e3
e7c42b83
00870713
01071a93
000ba503
010ada93
002a9593
899fb0ef
dc0504e3
00aba023
015b9223
8a0ff06f
000106b7
ff668693
dae6e8e3
e7c42783
00870713
0007a503
01071793
0107d793
00279593
e6f42823
85dfb0ef
d80506e3
e7c42703
e7042783
00a72023
00f71223
c2cff06f
e7042783
0007a703
00a70023
9cdff06f
e6e42223
984ff06f
e6e42223
b04ff06f
e6e42223
ad8ff06f
000b2503
815fb0ef
ce050ce3
00ab2023
cf1ff06f
017d0d33
8d551c63
e9042783
00400713
8ce78863
fff48493
8c8ff06f
e5042503
00371593
00070b13
fdcfb0ef
e4a42823
d00500e3
e5442703
001b1793
01250a33
00a72023
e4f42623
f1cff06f
0049a703
0009a683
5e975a63
0309a583
00000913
04098a13
00e686b3
00d9a023
00090a93
00048b13
00e90933
40e484b3
46058063
01458663
000c8513
fecef0ef
03c9a703
0209a823
00e9a223
44070263
0389a683
00000593
00d9a023
fa974ee3
015b0933
40970733
009686b3
00e9a223
00d9a023
012d0d33
e6442903
dd1fe06f
e7042783
e4042623
e4042823
e4f42223
e4042a23
e8440a13
d5cff06f
0009a683
0006c703
fc070793
00878733
f0074703
00071463
cb9fe06f
0049a703
00168693
00d9a023
fff70713
00e9a223
00100693
fad482e3
04098a13
02e05e63
0009a783
0007c703
fc070713
00870733
f0074703
f80702e3
0049a703
00178793
00190913
fff70713
00e9a223
00f9a023
f72484e3
fce046e3
0309a583
46058463
01458663
000c8513
f04ef0ef
03c9a783
0209a823
00f9a223
44078663
0389a783
00f9a023
fa1ff06f
00100593
c11ff06f
e4042c23
00000a93
00000a13
e8440b93
a6cff06f
e7042783
e4042c23
e4042a23
e4f42623
e6042823
00000913
e81fe06f
000a0913
00000b93
00000a13
919ff06f
ffe00793
b2f50263
000ba503
e5642823
ee1f60ef
e5042703
34051263
00300793
016d0d33
acfc1a63
e9042783
00400713
ace78663
fff48493
ac4ff06f
00294683
008aea93
00290913
b59fe06f
00294683
002aea93
00290913
b49fe06f
001b9b93
000a8513
000b8593
e5042c23
dc0fb0ef
00050a93
ae0502e3
e5842803
01250b33
00aa2023
8ddff06f
000b0a13
00000b93
00000b13
965ff06f
000a0b93
e7642823
e4042c23
00000a93
00000a13
990ff06f
e7042903
e4042c23
e4042a23
e6042823
dadfe06f
e5442a03
e4042623
e4042823
e4042a23
b94ff06f
ff010113
00f10793
ff07f793
e6f42e23
0007a023
0007a223
83cff06f
004af713
2a070863
01a69023
e6c42823
bbdfe06f
0309a583
36058e63
01058a63
000c8513
e5042c23
d80ef0ef
e5842803
03c9a783
0209a823
00f9a223
34078c63
0389a703
00e9a023
839ff06f
0009a683
0006c703
00ed8733
00074703
00877713
e8071463
0049a703
00168693
00d9a023
fff70713
00e9a223
00100693
00100a13
e6d48463
04098913
04e05063
0009a783
0007c703
00ed8733
00074703
00877713
e4071463
0049a703
00178793
001a0a13
fff70713
00e9a223
00f9a023
fd4496e3
014d0d33
e28ff06f
0309a583
24058e63
01258663
000c8513
cd0ef0ef
03c9a783
0209a823
00f9a223
24078063
0389a783
00f9a023
f9dff06f
e6042c23
a0dfe06f
00c9d703
0109a603
0009a223
02076713
00c9a023
00e99623
000b9463
d2dfe06f
931ff06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
b6090663
911ff06f
001af713
d6071e63
002afa93
d60a8a63
e6042783
00011737
b0870713
e7442683
00000613
000b0593
000c8513
20e78a63
ae1fd0ef
00050693
00058713
e7042783
0007a603
00d62023
00e62223
d40ff06f
00080b13
b0090863
e9840793
016787b3
fff7c583
fffb0b13
00098613
000c8513
d28fe0ef
fe0b12e3
aecff06f
00000b13
870ff06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
000c0b13
e5842c03
835a10e3
865ff06f
00c9d703
0109a683
e7142a23
02076713
0009a223
00d9a023
00e99623
b88ff06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
bc0916e3
825ff06f
0309a583
18058663
e5442783
00f58663
000c8513
b64ef0ef
03c9a783
0209a823
00f9a223
16078663
0389a783
00f9a023
fe5fe06f
e5042703
000b1463
ff1fe06f
00070493
e9840793
009787b3
fff7c583
fff48493
00098613
000c8513
c50fe0ef
fe0492e3
fc9fe06f
e7042483
0004a503
a98fb0ef
00051463
bc1fe06f
00a4a023
bb9fe06f
001af713
02071063
002afa93
000a8c63
41fd5713
01a6a023
00e6a223
e6c42823
8f9fe06f
01a6a023
e6c42823
8edfe06f
e5442483
00458593
0004a503
a48fb0ef
9e050063
00a4a023
9d8ff06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
addff06f
fff00793
e6f42c23
fe4fe06f
00c9d703
0109a683
0009a223
02076713
00d9a023
00e99623
014d0d33
ba8ff06f
000a8513
00369593
e4f42823
9e4fb0ef
00050a93
f0050463
e5042783
00aa2023
00f50bb3
e5842783
00179793
e4f42c23
ebdfe06f
00048913
a65ff06f
864fe0ef
00050693
00058713
df1ff06f
00c9d703
0109a683
415b0ab3
02076713
00d9a023
0009a223
00e99623
001a8593
015d0d33
000b0913
f1cff06f
00c9d703
0109a603
0009a223
02076713
00c9a023
00e99623
e60b1c63
e81fe06f
e7842783
e8078463
00c9d783
0407f793
e6079e63
e7c42783
f00fe06f
000a2b03
00fb0463
810ff06f
84cff06f
e1010113
1e112623
1f212023
1d812423
1da12023
00058c13
00060913
00d12a23
1e812423
1e912223
1d312e23
1d412c23
1d512a23
1d612823
1d712623
1d912223
1bb12e23
00050d13
d3cf90ef
00052783
00078513
02f12823
f64f00ef
00cc5783
0e012823
0e012a23
0e012c23
0e012e23
0807f793
02a12623
00078863
010c2783
00079463
3b80106f
10c10793
00078893
0ef12223
000247b7
47078793
00f12c23
000247b7
68478793
00090b13
00f12423
000b4783
0e012623
0e012423
02012023
02012a23
02012c23
02012e23
04012223
04012423
00012623
00088c93
22078263
000b0413
02500713
2ce78263
00144783
00140413
fe079ae3
416404b3
21640263
0ec12703
0e812783
016ca023
00970733
00178793
009ca223
0ee12623
0ef12423
00700713
008c8c93
28f74a63
00c12703
00044783
00970733
00e12623
1c078263
fff00313
00144483
0c0103a3
00140413
00000993
00000a13
05a00913
00900a93
02a00b93
00030d93
00140413
fe048793
04f96463
01812703
00279793
00e787b3
0007a783
00078067
00000993
fd048693
00044483
00299793
013787b3
00179793
00f689b3
fd048693
00140413
fedaf2e3
fe048793
fcf970e3
14048463
14910623
0c0103a3
00100a93
00100b93
14c10b13
00012823
00000313
02012423
02012223
00012e23
002a7f93
000f8463
002a8a93
084a7913
0ec12783
00091663
415986b3
40d040e3
0c714703
02070a63
0e812703
0c710693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
2ae6c863
020f8a63
0e812703
0c810693
00dca023
00278793
00200693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
4ce6c2e3
08000713
1ce900e3
41730db3
2bb042e3
100a7713
06071ee3
0e812703
017787b3
016ca023
00170713
017ca223
0ef12623
0ee12423
00700693
36e6cc63
008c8c93
004a7a13
000a0663
415984b3
38904263
0159d463
000a8993
00c12703
01370733
00e12623
300792e3
01012783
0e012423
00078863
01012583
000d0513
eb1ee0ef
10c10c93
00040b13
000b4783
de0792e3
0ec12783
00078463
2c90106f
00cc5783
0407f793
00078463
32c0206f
1ec12083
1e812403
00c12503
1e412483
1e012903
1dc12983
1d812a03
1d412a83
1d012b03
1cc12b83
1c812c03
1c412c83
1c012d03
1bc12d83
1f010113
00008067
000d0513
a24f90ef
00452783
00078513
04f12423
c4cf00ef
00050793
000d0513
00078493
04f12223
a00f90ef
00852783
02f12e23
00048463
7b10006f
00044483
dcdff06f
00044483
020a6a13
dc1ff06f
416404b3
d56418e3
00044783
d85ff06f
0e410613
000c0593
000d0513
364070ef
f40510e3
10c10c93
d59ff06f
008a7793
000d8313
740790e3
01412783
0b010513
01b12823
00778793
ff87f793
0047a603
0007a583
00878793
00f12a23
7710e0ef
0b012603
0b412683
0b812703
0bc12783
01012303
0f010513
00612823
0ef12e23
0ec12823
0ed12a23
0ee12c23
8ccf90ef
0ca12623
00200793
01012303
00f51463
4780106f
00100793
00f51463
5d80106f
06100793
00f49463
6190106f
04100793
00f49463
0380206f
fdf4f713
fff00793
02e12423
00f31463
1990106f
04700793
00f71463
1a40206f
0fc12d83
05412023
0f012e03
0f412e83
0f812f03
100a6793
000dd463
72d0106f
04012c23
00078a13
00012823
fbf48793
02500713
00f77463
6b40106f
00024737
00279793
5dc70713
00e787b3
0007a783
00078067
0e410613
000c0593
000d0513
04612623
05f12023
230070ef
0e0516e3
0ec12783
04c12303
04012f83
10c10c93
d29ff06f
0e812483
02012683
00100713
016ca023
00178793
00148493
008c8d93
3ad75ae3
00100713
00eca223
0ef12623
0e912423
00700713
50974ae3
02c12703
03012683
00148493
00e787b3
00eda223
00dda023
0ef12623
0e912423
00700713
008d8d93
509746e3
0f012703
0a010593
0b010513
0ae12823
0f412703
00f12e23
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
6290b0ef
02012783
fff78913
01c12783
360500e3
001b0813
00148493
012787b3
010da023
012da223
0ef12623
0e912423
00700713
008d8d93
30974ae3
03812683
0d410713
00148493
00f687b3
00eda023
00dda223
0ef12623
0e912423
00700713
008d8c93
c8975ae3
0e410613
000c0593
000d0513
100070ef
7a051e63
0ec12783
10c10c93
c75ff06f
01000693
0e812703
0096c463
6d10106f
000246b7
67468d93
01000913
00700a13
00c0006f
ff048493
04995663
01078793
00170713
01bca023
012ca223
0ef12623
0ee12423
008c8c93
fcea5ee3
0e410613
000c0593
000d0513
094070ef
74051863
ff048493
0ec12783
0e812703
10c10c93
fa994ee3
009787b3
00170713
01bca023
009ca223
0ef12623
0ee12423
00700693
bee6d8e3
0e410613
000c0593
000d0513
04c070ef
70051463
0ec12783
bd5ff06f
01412783
0c0103a3
0007ab03
00478913
000b1463
25c0106f
fff00793
54fd8ce3
000d8613
00000593
000b0513
01b12a23
be8f90ef
00a12823
01412303
00051463
4fd0106f
01012783
41678bb3
0c714783
fffbca93
41fada93
01212a23
00012823
02012423
02012223
00012e23
015bfab3
00000313
a80780e3
001a8a93
a79ff06f
01412703
0c0103a3
00100a93
00072783
00470713
00e12a23
14f10623
00100b93
14c10b13
a3dff06f
01412783
0007a983
00478793
3009dee3
413009b3
00f12a23
00044483
004a6a13
9b1ff06f
01412683
020a7793
00468713
32079ce3
010a7793
00078463
1700106f
040a7793
00078463
3580106f
200a7a13
000a1463
1580106f
01412783
00e12a23
00c12703
0007a783
00040b13
00e78023
af1ff06f
00044483
06c00793
3ef48ee3
010a6a13
94dff06f
01412703
ffff87b7
8307c793
0cf11423
00470793
000d8313
00f12a23
00072d83
000257b7
ea478793
02f12a23
00000913
002a6a93
00200793
07800493
00000693
0cd103a3
fff00693
1cd30863
012de6b3
f7fafa13
1c069063
22031663
04079ee3
001afb93
1b010b13
240b92e3
0c714783
00030a93
01735463
000b8a93
00012823
02012423
02012223
00012e23
ea079ee3
935ff06f
000d8313
010a6a13
020a7793
0c0788e3
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
bffa7a93
00000793
f75ff06f
00044483
06800793
2ef486e3
040a6a13
86dff06f
000d8313
010a6a93
020af793
0a078ae3
01412783
00778b13
ff8b7b13
008b0793
00f12a23
000b2d83
004b2903
00100793
f2dff06f
00044483
008a6a13
82dff06f
00044483
001a6a13
821ff06f
0c714783
00044483
80079ae3
02000793
0cf103a3
809ff06f
00044483
080a6a13
ffcff06f
00044483
00140713
01749463
6190106f
fd048693
00070413
00000d93
fedae063
00044483
002d9793
01b787b3
00179793
00d78db3
fd048693
00140413
fedaf2e3
fbcff06f
02b00793
00044483
0cf103a3
fa8ff06f
000d8313
010a6a13
020a7793
02078ee3
01412783
00778b13
ff8b7b13
004b2783
000b2d83
008b0713
00e12a23
00078913
0407c6e3
fff00793
000a0a93
00f30863
012de7b3
f7fa7a93
6c078263
48091ae3
00900793
49b7e6e3
030d8d93
1bb107a3
000a8a13
00100b93
1af10b13
e5dff06f
000a0a93
00100693
fcd78ae3
00200693
06d78c63
1b010b13
01d91713
007df793
003ddd93
03078793
01b76db3
00395913
fefb0fa3
012de733
000b0613
fffb0b13
fc071ce3
001af693
06068a63
03000693
06d78663
ffe60613
1b010793
fedb0fa3
40c78bb3
000a8a13
00060b13
dedff06f
00100713
00e79463
27d0106f
00200713
000a0a93
f8e798e3
03412683
1b010b13
00fdf793
00f687b3
0007c703
004ddd93
01c91793
01b7edb3
00495913
feeb0fa3
012de7b3
fffb0b13
fc079ce3
1b010793
41678bb3
000a8a13
d91ff06f
06500713
a0975ae3
0f012703
0a010593
0b010513
0ae12823
0f412703
04f12023
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
09d0b0ef
04012783
40051663
0e812703
000256b7
ed468693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
4ce6c6e3
0cc12703
02012683
70d75e63
03012703
02c12683
008c8c93
feecac23
0e812703
00d787b3
fedcae23
00170713
0ef12623
0ee12423
00700693
02e6cae3
02012703
fff70493
ee905463
01000693
0e812703
4896dce3
01000913
00700b93
00c0006f
ff048493
489952e3
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
311060ef
1c051663
0ec12783
0e812703
10c10c93
fb5ff06f
41598933
e5205063
01000613
0e812703
09265463
04812023
01000e13
000c0413
00700d93
00090c13
00030913
00c0006f
ff0c0c13
058e5a63
00812683
01078793
00170713
00dca023
01cca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
00040593
000d0513
291060ef
40051ee3
01000e13
ff0c0c13
0ec12783
0e812703
10c10c93
fb8e4ae3
00090313
000c0913
00040c13
04012403
00812683
012787b3
00170713
00dca023
012ca223
0ef12623
0ee12423
00700693
008c8c93
d8e6d463
0e410613
000c0593
000d0513
04612023
229060ef
0e051263
04012303
0ec12783
10c10c93
41730db3
d7b05263
01000613
0e812703
07b65463
01000313
00700913
00c0006f
ff0d8d93
05b35a63
00812683
01078793
00170713
00dca023
006ca223
0ef12623
0ee12423
008c8c93
fce95ce3
0e410613
000c0593
000d0513
1bd060ef
06051c63
01000313
ff0d8d93
0ec12783
0e812703
10c10c93
fbb34ae3
00812683
01b787b3
00170713
00dca023
01bca223
0ef12623
0ee12423
00700693
008c8c93
cce6d663
0e410613
000c0593
000d0513
169060ef
02051263
0ec12783
10c10c93
cacff06f
0e410613
000c0593
000d0513
149060ef
ce050863
01012583
d0058e63
000d0513
ba4ee0ef
d10ff06f
01000613
0e812703
00d64463
64c0106f
00024637
67460d93
05212623
04812823
000d8913
000d0413
000a8d93
01000e13
00098a93
00700293
00048993
05f12023
000c0493
00068d13
000b0c13
00030b13
00c0006f
ff0d0d13
05ae5a63
01078793
00170713
012ca023
01cca223
0ef12623
0ee12423
008c8c93
fce2dee3
0e410613
00048593
00040513
0a5060ef
1a051ae3
01000e13
ff0d0d13
0ec12783
0e812703
10c10c93
00700293
fbae4ae3
000d0693
000b0313
00040d13
000c0b13
04012f83
00048c13
05012403
00098493
000a8993
000d8a93
00090d93
04c12903
00d787b3
00170713
00dca223
01bca023
0ef12623
0ee12423
00700693
008c8c93
b0e6d463
0e410613
000c0593
000d0513
04612623
05f12023
019060ef
ec051ae3
0ec12783
04c12303
04012f83
10c10c93
ad8ff06f
0e410613
000c0593
000d0513
04612023
7ec060ef
ea0514e3
0ec12783
04012303
10c10c93
b1cff06f
0cc12603
00c05ae3
01c12703
02012683
00070493
3ee6ce63
02905663
0e812703
009787b3
016ca023
00170713
009ca223
0ef12623
0ee12423
00700693
008c8c93
34e6cee3
fff4c713
41f75713
00e4f4b3
01c12703
409704b3
4c904263
01c12683
400a7713
00db04b3
50071e63
0cc12683
02012703
00e6c663
001a7713
340704e3
03012703
02c12603
008c8c93
feecac23
0e812703
00c787b3
feccae23
00170713
0ef12623
0ee12423
00700613
00e65463
3f00106f
02012703
00eb0833
40d70633
40980933
01265463
00060913
03205863
0e812703
012787b3
009ca023
00170713
012ca223
0ef12623
0ee12423
00700693
008c8c93
00e6d463
4280106f
fff94713
41f75713
00e97933
412604b3
a4905663
01000693
0e812703
7e96de63
01000913
00700b93
00c0006f
ff048493
7e995463
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
674060ef
d20518e3
0ec12783
0e812703
10c10c93
fb5ff06f
940316e3
000a8a13
00000313
00000b93
1b010b13
fa8ff06f
001a7613
c4061663
00eca223
0ef12623
0e912423
00700713
ce975a63
0e410613
000c0593
000d0513
61c060ef
cc051ce3
0ec12783
0e812483
10c10d93
cd0ff06f
cd205663
01000713
052758e3
01000b93
00700b13
00c0006f
ff090913
032bdee3
00812703
01078793
00148493
00eda023
017da223
0ef12623
0e912423
008d8d93
fc9b5ce3
0e410613
000c0593
000d0513
5b4060ef
c60518e3
0ec12783
0e812483
10c10d93
fb5ff06f
01412703
010a7793
00072d83
00470713
00e12a23
14079a63
040a7793
14078263
010d9d93
010ddd93
00000913
f24ff06f
01412703
010af793
00072d83
00470713
00e12a23
02079663
040af793
00078c63
010d9d93
010ddd93
00000913
00100793
e6cff06f
200af793
00078463
0ffdfd93
00000913
00100793
e54ff06f
01412703
010a7793
00072d83
00470713
00e12a23
0c079263
040a7793
0a078a63
010d9d93
410ddd93
41fdd913
00090793
fa07de63
01b037b3
41200933
40f90933
41b00db3
000a0a93
02d00693
00100793
e04ff06f
0e410613
000c0593
000d0513
4c0060ef
b6051ee3
0ec12783
0e812483
10c10d93
ad0ff06f
0e410613
000c0593
000d0513
49c060ef
b4051ce3
0ec12783
0e812483
10c10d93
ad8ff06f
001a7713
00071463
800ff06f
8ddff06f
000d8313
f10ff06f
00044483
00f12a23
ea1fe06f
03000793
1af107a3
1af10b13
db4ff06f
200a7793
080790e3
41fdd913
00090793
f08ff06f
200a7793
080790e3
00000913
de4ff06f
00c12603
0006a783
00e12a23
41f65693
00c7a023
00d7a223
00040b13
fddfe06f
01412703
00072783
00470713
00e12a23
0007a603
0047a683
0087a703
00c7a783
8e0ff06f
03c12783
00044483
00079463
e19fe06f
0007c783
00079463
e0dfe06f
400a6a13
e05fe06f
00068493
c09044e3
c2dff06f
000d8313
000a0a93
d8cff06f
000257b7
ea478793
000d8313
02f12a23
020a7793
2a078863
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
001a7793
00078e63
012de7b3
00078a63
03000793
0cf10423
0c9104a3
002a6a13
bffa7a93
00200793
c80ff06f
00144483
200a6a13
00140413
d7dfe06f
0e410613
000c0593
000d0513
330060ef
9e0516e3
0ec12783
10c10c93
fb4ff06f
00144483
020a6a13
00140413
d4dfe06f
000257b7
eb878793
000d8313
02f12a23
f61ff06f
000d8313
c84ff06f
04000593
000d0513
a70ee0ef
00ac2023
00ac2823
00051463
3700106f
04000793
00fc2a23
c29fe06f
000b0513
b54ef0ef
00050b93
accff06f
01000693
0e812703
5c96dc63
01000b93
00700d93
00c0006f
ff048493
5c9bd263
00812683
01078793
00170713
00dca023
017ca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
000c0593
000d0513
268060ef
920512e3
0ec12783
0e812703
10c10c93
fb5ff06f
02012703
02412b83
00812e23
00eb0733
05412023
05312623
03512223
02812983
03612423
03c12403
04412a03
04812a83
00700d93
01000913
000c8693
00070b13
080b8663
08099663
fff40413
fffb8b93
0e812703
014787b3
0156a023
00170713
0146a223
0ef12623
0ee12423
00868693
12edcc63
00044603
409b0cb3
01965463
00060c93
03905663
0e812603
019787b3
0096a023
00160613
0196a223
0ef12623
0ec12423
30cdcc63
00044603
00868693
fffcc513
41f55513
00acf733
40e60cb3
01904c63
00c484b3
f60b9ee3
3c0988e3
fff98993
f7dff06f
0e812603
01994863
0580006f
ff0c8c93
05995863
00812703
01078793
00160613
00e6a023
0126a223
0ef12623
0ec12423
00868693
fccddce3
0e410613
000c0593
000d0513
134060ef
fe051863
ff0c8c93
0ec12783
0e812603
10c10693
fb994ce3
00812703
019787b3
00160613
00e6a023
0196a223
0ef12623
0ec12423
42cdc0e3
00044603
00868693
00c484b3
f65ff06f
01412703
010a7793
00072d83
00470713
00e12a23
02079263
040a7793
00078a63
010d9d93
010ddd93
00000913
d45ff06f
200a7793
4c079e63
00000913
d35ff06f
0e410613
000c0593
000d0513
09c060ef
f4051c63
0ec12783
10c10693
eb1ff06f
1b010b13
00000793
00812823
00912e23
000b0413
03312223
000c0b13
000d8493
00090993
03c12d83
400afa13
0ff00b93
00030c13
00078913
0240006f
00a00613
00000693
00048513
00098593
469070ef
3e098463
00050493
00058993
00a00613
00000693
00048513
00098593
208080ef
03050513
fea40fa3
00190913
fff40413
fa0a0ee3
000dc683
fad91ae3
fb7908e3
36099463
00900793
3697e063
000c0313
1b010793
000b0c13
00040b13
01c12483
02412983
01012403
03b12e23
03212023
41678bb3
000a8a13
920ff06f
0e812703
000256b7
ed468693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
06e6ce63
1e061863
02012683
001a7713
00d76733
00071463
af9fe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
60e6c263
02012683
00170713
0168a023
00f687b3
00d8a223
0ef12623
0ee12423
00700693
00888c93
00e6c463
a9dfe06f
e09fe06f
0e410613
000c0593
000d0513
705050ef
dc051063
0cc12603
0ec12783
10c10c93
f69ff06f
00040d13
00048c13
da4ff06f
0e410613
000c0593
000d0513
6d5050ef
d8051863
0ec12783
10c10c93
b1cff06f
00812683
009787b3
009ca223
00dca023
00170713
0ef12623
0ee12423
00700693
00e6c463
a1dfe06f
d8dfe06f
0e410613
000c0593
000d0513
689050ef
d4051263
00044603
0ec12783
10c10693
cd5ff06f
00040c13
d2cff06f
0f012783
0a010593
0b010513
0af12823
0f412783
0a012023
0a012223
0af12a23
0f812783
0a012423
0a012623
0af12c23
0fc12783
0af12e23
4f50a0ef
320540e3
0c714783
04700713
1c975e63
00025837
e9880b13
00012823
02012423
02012223
00012e23
f7fa7a13
00300a93
00300b93
00000313
00078463
e2dfe06f
8a5fe06f
01412783
00040b13
0007a783
00e12a23
00c12703
00e7a023
99dfe06f
00600793
000d8b93
1bb7e663
00025837
000b8a93
01212a23
ecc80b13
855fe06f
00812703
012787b3
00148493
00eda023
c4dfe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
42e6c663
e20654e3
ff000693
40c004b3
3ed658e3
01000913
00700b93
00c0006f
ff048493
3c995ee3
00812683
01078793
00170713
00d8a023
0128a223
0ef12623
0ee12423
00888893
fcebdce3
0e410613
000c0593
000d0513
515050ef
bc051863
0ec12783
0e812703
10c10893
fb5ff06f
0fc12783
3a07d863
02d00793
0cf103a3
04700713
229750e3
00025837
ea080b13
ec9ff06f
00812683
009787b3
00170713
00dca023
009ca223
0ef12623
0ee12423
00700693
008c8c93
d2e6de63
0e410613
000c0593
000d0513
4a5050ef
b6051063
0ec12783
10c10c93
d1cff06f
04412783
04812583
00000913
40f40433
00078613
00040513
8d4fa0ef
001dc583
00a00613
00000693
00b03833
00048513
00098593
010d8db3
085070ef
c21ff06f
00900793
c097ece3
c5dff06f
00025837
e9480b13
e29ff06f
0e410613
000c0593
000d0513
42d050ef
ae051463
0ec12783
10c10c93
c8cff06f
00600b93
e55ff06f
02012703
00eb0833
40d70633
40980933
d3265463
00060913
d20ff06f
01412783
00e12a23
00c12703
0007a783
00040b13
00e79023
fa8fe06f
0ffdfd93
00000913
859ff06f
018d9d93
418ddd93
41fdd913
00090793
e85fe06f
0ffdfd93
00000913
d65fe06f
00030693
00200613
0b010a93
0d010793
0cc10713
0dc10813
000a8593
000d0513
04612823
04d12623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
0bb12e23
ea8f60ef
02812703
04700793
01c12f03
02012e83
02412e03
04c12683
05012303
00050b13
64f70863
04600793
00d50933
06f71ee3
00054703
03000793
2ef700e3
0a010b93
0cc12783
00f90933
000b8593
000a8513
00612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
0a012023
0a012223
0a012423
0a012623
7a40a0ef
01c12303
00090693
02050263
0dc12683
0126fe63
03000713
00168793
0cf12e23
00e68023
0dc12683
ff26e8e3
416687b3
02f12023
0cc12703
04700793
00e12e23
02812703
52f70463
02812703
04600793
02f700e3
01c12783
02812603
04100693
fff78b93
0d712623
0ff4f793
00000713
00d61863
00f78793
0ff7f793
00100713
0cf10a23
02b00793
000bda63
01c12783
00100b93
40fb8bb3
02d00793
0cf10aa3
00900793
0b77d6e3
0e310a13
000a0913
00a00593
000b8513
c0dec0ef
03050793
fef90fa3
000b8513
00a00593
b75ec0ef
000b8a93
06300793
00090d93
00050b93
fff90913
fd57c6e3
03050693
0ff6f693
ffed8793
fed90fa3
2947f0e3
0d610713
0080006f
0007c683
00d70023
00178793
00170713
ff4798e3
0e510793
0d610713
41b787b3
00f707b3
0d410713
40e787b3
02f12c23
02012703
03812683
00100793
00d70bb3
0ce7d6e3
02c12783
00fb8bb3
04012783
fffbca93
41fada93
bff7fa13
100a6a13
015bfab3
02012423
02012223
00012e23
05812783
40078a63
02d00793
0cf103a3
00000313
001a8a93
c18fe06f
0e410613
000c0593
000d0513
151050ef
d2cfe06f
0c714783
c59ff06f
0e410613
000c0593
000d0513
135050ef
00050463
fedfe06f
0cc12603
0ec12783
0e812703
10c10893
9c065ce3
bb1ff06f
00600313
e74fe06f
00130693
00200613
d5dff06f
00030693
00300613
d51ff06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
09d0d0ef
0cc10613
ae5f90ef
00058613
00050593
000a8513
5080d0ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
0710a0ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
4d00a0ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000257b7
eb878793
02f12223
fff30913
06912023
07312423
07912823
07a12a23
07812c23
01c12483
00090c13
04812e23
07412223
06612623
000b0c93
07612e23
00068d13
000e0d93
000e8913
000f0993
0480006f
000b8593
000a8513
02c12023
01f12e23
0bf12c23
0ac12e23
0b612823
0b412a23
0a012023
0a012223
0a012423
0a012623
4280a0ef
fffc0c13
00090f93
00098613
0e050263
400307b7
00048613
000b8593
000a8513
08f12e23
0ba12023
0bb12223
0b212423
0b312623
08012823
08012a23
08012c23
7380a0ef
000a8513
0100d0ef
00050593
00050413
000a8513
0b012a03
0b412983
0b812b03
0bc12903
1040d0ef
0b012683
04c12603
00048593
08d12023
0b412683
000b8513
09412823
08d12223
0b812683
09312a23
09612c23
08d12423
0bc12683
09212e23
08d12623
2950b0ef
02412783
0a012b03
0a412a03
008786b3
0006c683
0a812f83
0ac12603
05912a23
00dc8023
05812823
fff00793
001c8c93
000b0d13
000a0d93
000f8913
00060993
eefc10e3
06c12303
000b0393
000a0293
3ffe0937
000b8593
000a8513
02612023
00812e23
06012483
05c12403
06412a03
0a712823
06712223
0a512a23
06512023
0bf12c23
05f12e23
0ac12e23
04c12623
0a012023
0a012223
0a012423
0b212623
3a40a0ef
000c8d93
06812983
07012c83
07412d03
07812c03
07c12b03
02012303
40a04463
000b8593
000a8513
2ac0a0ef
02012303
00051863
01c12783
0017f913
3e091463
05012783
03000693
00178713
00ed8733
0007c863
001d8d93
fedd8fa3
ffb71ce3
416d87b3
02f12023
b01ff06f
02812b03
02012703
02812e23
04012a03
00eb0733
01c12403
04c12983
02412a83
00068c93
00976463
e25fe06f
00070493
e1dfe06f
01c12703
ffd00793
00f74463
02e35463
ffe48493
fdf4f793
02f12423
acdff06f
0c714783
00000313
00078463
d90fe06f
808fe06f
02012783
01c12703
30f74263
04012783
01c12703
0017f793
00070b93
00078663
02c12783
00f70bb3
04012783
4007f793
00078663
01c12783
44f04463
fffbca93
41fada93
015bfab3
06700493
02012423
02012223
b81ff06f
04012783
00d50933
0017f793
22079663
0dc12683
a21ff06f
0e410613
000c0593
000d0513
4d0050ef
00050463
b89fe06f
00044603
0ec12783
10c10693
00c484b3
b2cff06f
07800793
03000713
0ce10423
002a6713
0cf104a3
04e12023
06300793
00012823
14c10b13
3667c863
0fc12d83
fdf4f793
02f12423
04012c23
0f012e03
0f412e83
0f812f03
102a6a13
120dc063
06100793
00f48463
9f0fe06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
4040d0ef
0cc10613
e4cf90ef
00058613
00050593
000a8513
0700d0ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
3d80a0ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
0380a0ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000257b7
ea478793
02f12223
b69ff06f
00012823
00078a13
800007b7
01b7cdb3
02d00793
04f12c23
ed5ff06f
0e410613
000c0593
000d0513
328050ef
00050463
9e1fe06f
0cc12683
0ec12783
10c10c93
bf1fe06f
02d00793
0cf103a3
ce0ff06f
0c714783
01212a23
02012423
02012223
00012e23
00030a93
00030b93
00000313
00078463
b18fe06f
d91fd06f
00024637
67460d93
a7dfe06f
00025837
e9c80b13
cacff06f
0a010b93
f9cff06f
0e410613
000c0593
000d0513
2a8050ef
00050463
961fe06f
0cc12483
02012703
0ec12783
10c10c93
40970633
bb1fe06f
05800793
dd5ff06f
04012783
01c12703
0017f793
0067e7b3
2ae05063
28079463
01c12b83
06600493
04012783
4007f793
18079663
fffbca93
41fada93
015bfab3
d45ff06f
02012783
02c12703
06700493
00e78bb3
01c12783
fcf048e3
40fb8bb3
001b8b93
fffbca93
41fada93
015bfab3
d15ff06f
000246b7
67468d93
990fe06f
000a0a93
cf0fe06f
05412783
000d8713
0cf12e23
02412783
fffdc683
00f7c603
02d61063
03000593
feb70fa3
0dc12703
fff70793
0cf12e23
fff74683
fed606e3
00168613
03900593
0ff67613
00b68663
fec70fa3
bf1ff06f
02412783
00a7c603
fec70fa3
be1ff06f
0d610793
00071863
03000793
0cf10b23
0d710793
1b010713
030b8b93
40e78733
01778023
0dd70793
02f12c23
fb8ff06f
00812683
009787b3
00170713
00d8a023
0098a223
0ef12623
0ee12423
00700693
00888893
a0e6d463
0e410613
000c0593
000d0513
138050ef
00050463
ff0fe06f
0ec12783
0e812703
10c10893
9e0ff06f
00130593
000d0513
00612823
898ed0ef
01012303
00050b13
1a050e63
00a12823
c75ff06f
00030463
e5dfd06f
00100313
e55fd06f
fff00793
00f12623
cd1fd06f
04012783
0017f793
f2078c63
f2cff06f
06700493
03c12603
0ff00713
00064783
16e78463
01c12683
00000513
00000593
00d7de63
40f686b3
00164783
04078463
00158593
00160613
fee794e3
02c12e23
00d12e23
02b12223
02a12423
02812783
02412703
04412583
00e78533
9a0ec0ef
01750bb3
fffbca93
41fada93
015bfab3
ee4ff06f
00064783
00150513
fbdff06f
0a010b93
000b8593
000a8513
04612623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
04d12823
0bb12e23
0a012023
0a012223
0a012423
0a012623
4c1090ef
01c12f03
02012e83
02412e03
04c12303
cc050a63
05012683
00100793
40d787b3
0cf12623
cc4ff06f
02c12783
06600493
00f70bb3
006b8bb3
d75ff06f
00079a63
00100a93
06600493
00100b93
abdff06f
02c12783
06600493
00178b93
006b8bb3
fffbca93
41fada93
015bfab3
a9dff06f
01412783
0007ad83
00478793
000dd463
fff00d93
00144483
00f12a23
00070413
9b5fd06f
00200793
02f12c23
db4ff06f
00c00793
00fd2023
fff00793
00f12623
b49fd06f
02012423
02012223
ecdff06f
00cc5783
0407e793
00fc1623
b1dfd06f
fe010113
00812c23
00058413
0305a583
00112e23
00912a23
01212823
01312623
01412423
04040793
06f58063
03442903
00191993
00098613
919f80ef
00050493
0a050463
01250a33
00050593
00090613
000a0513
b88f70ef
00000513
01442023
02942823
03342a23
01c12083
01812403
01412483
01012903
00c12983
00812a03
02010113
00008067
40000593
e35ec0ef
00050793
04050a63
04244703
40000693
02a42823
02d42a23
3ee50fa3
04144683
3fd50713
00000513
3ed78f23
04044683
3ed78ea3
01c12083
00e42023
01812403
01412483
01012903
00c12983
00812a03
02010113
00008067
fff00513
f7dff06f
fe010113
00112e23
00812c23
00912a23
01212823
01312623
fff00793
0ef58263
00058493
00050913
00060413
00050663
03852783
0c078a63
00c41783
01279713
02074463
06442703
000026b7
00d7e7b3
ffffe6b7
fff68693
00d77733
01079793
4107d793
06e42223
fdf7f793
01079713
00f41623
0047f693
01075713
00069e63
01077693
06068e63
00877713
0e071a63
0047e793
00f41623
03042703
0ff4f993
00442783
0ff4f493
06070a63
03442703
04e7d063
00042783
fff78713
00e42023
ff378fa3
00442783
00178793
00f42223
01c12083
01812403
01012903
00c12983
00048513
01412483
02010113
00008067
00040593
00090513
e19ff0ef
fa050ce3
fff00493
fcdff06f
e28ec0ef
00c41783
01279713
f4074ae3
f2dff06f
01042683
00042703
00068863
00e6f663
fff74683
06968a63
02f42e23
00300793
05340123
02f42a23
04040613
04240693
00100793
01c12083
02e42c23
02c42823
00d42023
00f42223
01812403
01012903
00c12983
00048513
01412483
02010113
00008067
00040593
00090513
960ec0ef
f6051ae3
00c41783
00042423
00042c23
ff77f793
ef1ff06f
fff70713
00178793
00e42023
00f42223
f1dff06f
04001737
00050793
9e472503
00058613
00078593
e35ff06f
0645a703
fd010113
000027b7
01612823
02112623
02812423
02912223
03212023
01312e23
01412c23
01512a23
01712623
01812423
00e7f7b3
00060b13
0a078863
00862783
00062b83
00058913
00050993
fff00a93
08078863
004bac03
000ba403
002c5a13
060a0663
00000493
00c0006f
00440413
049a0c63
00042583
00090613
00098513
738010ef
00148493
ff5512e3
fff00513
02c12083
02812403
000b2423
000b2223
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
008b2783
ffcc7c13
418787b3
00fb2423
008b8b93
f6079ce3
00000513
fadff06f
995f30ef
fa5ff06f
00862703
00070463
f05ff06f
00062223
00000513
00008067
ed010113
11312e23
11512a23
11712623
12112623
12812423
12912223
13212023
11412c23
11612823
11812423
11912223
11a12023
0fb12e23
00d12823
00050a93
00058993
00060b93
00050663
03852783
62078663
00c99703
000026b7
01071793
0107d793
00d7f633
02061863
0649a603
00d767b3
01079793
ffffe737
4107d793
fff70713
00e67733
00f99623
01079793
06e9a223
0107d793
0087f713
3e070a63
0109a703
3e070663
01a7f793
00a00713
40e78063
000247b7
69478793
00025b37
04c10493
00f12a23
00025937
800b0793
000b8c13
04912023
04012423
04012223
00012c23
00012e23
02012223
02012023
00012623
00f12423
81090913
00048b93
000c4783
26078263
000c0413
02500713
46e78263
00144783
00140413
fe079ae3
41840cb3
25840263
04812703
04412783
018ba023
00ec8733
00178793
019ba223
04e12423
04f12223
00700693
008b8b93
02f6d063
420700e3
04010613
00098593
000a8513
d91ff0ef
20051463
00048b93
00c12703
00044783
01970733
00e12623
1e078463
00144683
00140c13
02010da3
fff00a13
00012223
00000b13
05a00c93
00900d13
02a00613
001c0c13
fe068793
04fce863
01412703
00279793
00e787b3
0007a783
00078067
00012223
fd068793
00412583
000c4683
001c0c13
00259713
00b70733
00171713
00e787b3
00f12223
fd068793
fcfd7ee3
fe068793
fafcfce3
16068463
08d10623
02010da3
00100c93
00100d13
08c10413
00000a13
002b7f93
000f8463
002c8c93
04412703
084b7f13
04812783
00170693
00068613
000f1863
00412583
41958db3
0fb04ce3
03b14683
02068a63
03b10713
00178793
00eba023
00100713
00eba223
04f12423
04c12223
00700713
04c748e3
00060713
008b8b93
00160613
040f8c63
03c10713
00278793
00eba023
00200713
00eba223
04f12423
04c12223
00700713
08c750e3
32078ce3
04010613
00098593
000a8513
03e12423
c35ff0ef
0a051663
04412703
04812783
02812f03
00048b93
00170613
08000693
62df0a63
41aa0a33
71404263
00fd07b3
008ba023
01aba223
04f12423
04c12223
00700713
60c75463
12078ee3
04010613
00098593
000a8513
bddff0ef
04051a63
04812783
00048b93
004b7e13
000e0863
00412703
41970d33
13a044e3
00412403
01945463
000c8413
00c12703
00870733
00e12623
74079463
000c4783
04012223
00048b93
da0792e3
04812783
5e079ae3
00c9d783
0407f793
620792e3
12c12083
12812403
00c12503
12412483
12012903
11c12983
11812a03
11412a83
11012b03
10c12b83
10812c03
10412c83
10012d03
0fc12d83
13010113
00008067
000a8513
e04f60ef
00452783
00078513
02f12023
82ded0ef
00050793
000a8513
00078413
02f12223
de0f60ef
00852783
02a00613
00f12e23
320416e3
000c4683
dadff06f
000c4683
020b6b13
da1ff06f
010b6b13
020b7793
1a078063
01012783
00778793
ff87f793
0047a683
0007ad03
00878793
00f12823
00068c93
1a06c863
fff00693
000b0d93
00da0863
019d66b3
f7fb7d93
120688e3
1a0c9ae3
00900693
1ba6e6e3
030d0793
0ef107a3
000d8b13
00100d13
0ef10413
000a0c93
01aa5463
000d0c93
03b14783
00f037b3
00fc8cb3
d91ff06f
00098593
000a8513
878f30ef
500510e3
00c9d783
00a00713
01a7f793
c0e794e3
00e99783
c007c0e3
12812403
01012683
12c12083
12412483
12012903
11812a03
11012b03
10812c03
10412c83
10012d03
0fc12d83
000b8613
00098593
10c12b83
11c12983
000a8513
11412a83
13010113
4e90006f
010b6b13
020b7793
06078c63
01012783
00778793
ff87f793
0007ad03
0047ac83
00878793
00f12823
bffb7d93
00000693
00000613
02c10da3
fff00613
0cca0863
019d6633
f7fdfb13
5e061663
340a1463
02069ae3
001dfd13
0f010413
f00d0ae3
03000793
0ef107a3
0ef10413
f05ff06f
41840cb3
bb8418e3
00044783
c01ff06f
01012683
010b7713
0006a783
00468693
00d12823
14071e63
040b7713
14070663
01079d13
010d5d13
00000c93
f7dff06f
01012683
010b7713
0006a783
00468693
00d12823
14071063
040b7713
12070863
01079d13
410d5d13
41fd5c93
000c8693
e406dce3
02d00613
01a036b3
41900733
02c10da3
fff00613
40d70cb3
41a00d33
000b0d93
00100693
f2ca1ce3
00100613
e4c680e3
00200613
28c68863
0f010413
01dc9793
007d7693
003d5d13
03068693
01a7ed33
003cdc93
fed40fa3
019d67b3
00040593
fff40413
fc079ce3
001df793
28078663
03000793
28f68263
ffe58593
fef40fa3
0f010793
40b78d33
000d8b13
00058413
dfdff06f
dd9eb0ef
9d5ff06f
01012783
02010da3
0007a403
00478d93
20040ce3
fff00793
16fa02e3
000a0613
00000593
00040513
89df60ef
2c0502e3
40850d33
01b12823
00000a13
db5ff06f
01012703
02010da3
00100c93
00072783
00470713
00e12823
08f10623
00100d13
08c10413
b31ff06f
200b7713
24071ae3
00078d13
00000c93
e31ff06f
200b7713
220710e3
41f7dc93
00078d13
000c8693
d25ff06f
01012783
0007a703
00478793
00e12223
78075463
00412703
00f12823
40e00733
00e12223
000c4683
004b6b13
a65ff06f
000c4683
06c00793
12f68ae3
010b6b13
a51ff06f
000c4683
06800793
10f688e3
040b6b13
a3dff06f
010b6d93
020df793
62078063
01012783
00100693
00778793
ff87f793
0007ad03
0047ac83
00878793
00f12823
d99ff06f
000c4683
001b6b13
a01ff06f
03b14783
000c4683
9e079ae3
02000793
02f10da3
9e9ff06f
000c4683
080b6b13
9ddff06f
000c4683
001c0713
1cc688e3
fd068793
00070c13
00000a13
9cfd62e3
000c4683
002a1713
01470a33
001a1a13
00fa0a33
fd068793
001c0c13
fefd72e3
9a1ff06f
02b00793
000c4683
02f10da3
98dff06f
01012783
ffff86b7
8306c693
0007ad03
00478793
00f12823
000257b7
ea478793
02d11e23
00000c93
002b6d93
00f12c23
00200693
ce1ff06f
01012683
020b7793
00468713
6a079063
010b7793
020794e3
040b7793
08079ce3
200b7e13
000e0ce3
01012783
00e12823
00c12703
0007a783
00e78023
86dff06f
00100613
0ec68ce3
00200613
000b0d93
d6c69ce3
01812683
0f010413
00fd7793
00f687b3
0007c703
004d5d13
01cc9793
01a7ed33
004cdc93
fee40fa3
019d67b3
fff40413
fc079ce3
0f010793
40878d33
000d8b13
b89ff06f
00100713
000d0793
04812623
05a12823
05a12423
04e12223
00048b93
008b8b93
a19ff06f
00412683
41968db3
9db054e3
01000693
07b6dc63
01000e93
00700f13
0180006f
00270613
008b8b93
00068713
ff0d8d93
05bedc63
01078793
00170693
012ba023
01dba223
04f12423
04d12223
fcdf5ae3
14078863
04010613
00098593
000a8513
d80ff0ef
9e051ce3
04412703
01000e93
ff0d8d93
04812783
00048b93
00170613
00700f13
fbbec8e3
01b787b3
012ba023
01bba223
04f12423
04c12223
00700713
00060593
52c75e63
70078e63
04010613
00098593
000a8513
d28ff0ef
9a0510e3
04412703
41aa0a33
04812783
00048b93
00170613
914052e3
01000693
0746da63
01000893
00700d93
0180006f
00270613
008b8b93
00068713
ff0a0a13
0548da63
01078793
00170693
012ba023
011ba223
04f12423
04d12223
fcdddae3
04078e63
04010613
00098593
000a8513
cb4ff0ef
920516e3
04412703
01000893
ff0a0a13
04812783
00048b93
00170613
fb48cae3
014787b3
012ba023
014ba223
04f12423
04c12223
00700713
2cc74663
008b8b93
00160613
865ff06f
00100613
00000713
00048b93
f75ff06f
04010613
00098593
000a8513
c4cff0ef
8a0506e3
8c1ff06f
00100613
00000713
00048b93
e81ff06f
32078863
04010613
00098593
000a8513
03e12623
03f12423
c18ff0ef
880518e3
04412703
04812783
02c12f03
02812f83
00048b93
00170613
f88ff06f
3a079e63
03b14703
5e071463
2e0f8663
03c10793
04f12623
00200793
04f12823
00100613
00048b93
00060713
008b8b93
00170613
fa8ff06f
000b0d93
ad5ff06f
01000613
65b65063
000b8613
01000e93
00040b93
00700293
00098413
03f12423
000d8993
000c0d93
000a0c13
000f0a13
01c0006f
00270513
00860613
00068713
ff098993
053ede63
00170693
00812583
01078793
01d62223
00b62023
04f12423
04d12223
fcd2d8e3
08078663
04010613
00040593
000a8513
b3cff0ef
4a051863
04412703
01000e93
ff098993
04812783
00048613
00170513
00700293
fb3ec6e3
02812f83
000a0f13
00050593
000c0a13
000d8c13
00098d93
00040993
000b8413
00060b93
00812703
01b787b3
01bba223
00eba023
04f12423
04b12223
00700713
eeb740e3
008b8b93
00158613
00058713
e1cff06f
00000713
00100513
00048613
f41ff06f
04012223
004b7e13
0e0e0063
00412703
41970d33
0da05a63
00048b93
01000713
04412683
53a75263
01000d93
00700413
0180006f
00268613
008b8b93
00070693
ff0d0d13
05adda63
00812603
01078793
00168713
00cba023
01bba223
04f12423
04e12223
fce458e3
06078863
04010613
00098593
000a8513
a38ff0ef
ea051863
04412683
ff0d0d13
04812783
00048b93
00168613
fbadcae3
00812703
01a787b3
01aba223
00eba023
04f12423
04c12223
00700713
e4c75263
02078863
04010613
00098593
000a8513
9e8ff0ef
e6051063
04812783
e24ff06f
00100613
00000693
00048b93
f5dff06f
00412403
01945463
000c8413
00c12783
008787b3
00f12623
e14ff06f
ba0784e3
04010613
00098593
000a8513
99cff0ef
e0051a63
04412603
04812783
00048b93
00160613
d7cff06f
04012223
00048b93
bf4ff06f
ee0a1063
000d8b13
00000a13
00000d13
0f010413
ee0ff06f
01012683
010df713
0006a783
00468693
00d12823
02071463
040df713
00070c63
01079d13
010d5d13
00000c93
00100693
f6cff06f
200df713
38071063
00078d13
00000c93
00100693
f54ff06f
00100613
00000713
00048b93
cecff06f
140f9463
00000713
00100613
00048b93
cd8ff06f
400df793
03412423
03312623
000c8a13
000d0993
00000b13
01c12d03
0f010413
00078c93
0240006f
00a00613
00000693
00098513
000a0593
159050ef
280a0463
00050993
00058a13
00a00613
00000693
00098513
000a0593
6f9050ef
03050513
fea40fa3
001b0b13
fff40413
fa0c8ee3
000d4683
fb669ae3
0ff00793
fafb06e3
180a1863
00900793
1937e463
0f010793
01a12e23
02812a03
02c12983
40878d33
000d8b13
dc8ff06f
000c4683
00f12823
af0ff06f
04010613
00098593
000a8513
03e12623
03f12423
824ff0ef
c8051e63
04412703
04812783
02c12f03
02812f83
00048b93
00170613
b5cff06f
008b8b93
00160613
00058713
be4ff06f
00c12603
0006a783
00e12823
41f65693
00c7a023
00d7a223
9e4ff06f
01c12783
000c4683
a8078063
0007c783
a6078c63
400b6b13
a70ff06f
03c10793
04f12623
00200793
04f12823
00100713
00048b93
bd9ff06f
000b0d93
819ff06f
000257b7
ea478793
00f12c23
020b7793
06078063
01012783
00778793
ff87f793
0007ad03
0047ac83
00878793
00f12823
001b7613
00060e63
019d6633
00060a63
03000613
02c10e23
02d10ea3
002b6b13
bffb7d93
00200693
d7cff06f
000257b7
eb878793
00f12c23
020b7793
fa0794e3
01012603
010b7713
00062783
00460613
00c12823
06071e63
040b7713
06070663
01079d13
010d5d13
00000c93
f95ff06f
00040513
bf9ec0ef
00050d13
01b12823
00000a13
c60ff06f
02412783
02012583
00000b13
40f40433
00078613
00040513
f99f70ef
001d4583
00a00613
00000693
00b03733
00098513
000a0593
00ed0d33
748050ef
df5ff06f
200b7713
0c071e63
00078d13
00000c93
f29ff06f
00040993
b00ff06f
001c4683
200b6b13
001c0c13
928ff06f
001c4683
020b6b13
001c0c13
918ff06f
01012783
0007a783
00e12823
00c12703
00e7a023
858ff06f
00600793
000a0d13
0347ea63
00025337
000d0c93
01b12823
ecc30413
950ff06f
00900793
d737ece3
dc1ff06f
00100613
00000713
00048b93
a00ff06f
00600d13
fcdff06f
03b10793
04f12623
00100793
04f12823
00100613
00048b93
970ff06f
01012783
00e12823
00c12703
0007a783
00e79023
fe1fe06f
01879d13
418d5d13
41fd5c93
000c8693
b04ff06f
0ff7fd13
00000c93
e51ff06f
0ff7fd13
00000c93
be0ff06f
0ff7fd13
00000c93
00100693
bd8ff06f
04010613
00098593
000a8513
d89fe0ef
a00ff06f
000a0d13
01b12823
00000a13
af4ff06f
00068593
a7dff06f
00168613
b4dff06f
000b0d93
ac8ff06f
fff00793
00f12623
9d8ff06f
01012783
0007aa03
00478793
000a5463
fff00a13
001c4683
00f12823
00070c13
fe1fe06f
04001737
00050793
9e472503
00060693
00058613
00078593
e1dfe06f
00c5d783
0645ae03
00e5d303
01c5a883
0245a803
b8010113
ffd7f793
40000713
46812c23
00f11a23
00058413
07010793
00810593
46912a23
47212823
46112e23
00050913
07c12623
00611b23
03112223
03012623
00f12423
00f12c23
00e12823
00e12e23
02012023
db1fe0ef
00050493
02055c63
01415783
0407f793
00078863
00c45783
0407e793
00f41623
47c12083
47812403
47012903
00048513
47412483
48010113
00008067
00810593
00090513
d75ea0ef
fc0500e3
fff00493
fb9ff06f
040017b7
9307a783
00078067
02058463
0ff00793
00c7e863
00c58023
00100513
00008067
08a00793
00f52023
fff00513
00008067
00000513
00008067
040017b7
9e47a703
ff010113
00068793
00060813
00112623
00c72883
00050693
00058713
00078613
02080063
000257b7
fdc78793
000255b7
fec58593
00088513
210000ef
399040ef
00025837
e3c80793
e3c80813
fe1ff06f
ff010113
00060693
00000613
00112623
f99ff0ef
00050593
00000693
00000613
00000513
3790406f
fe010113
00812c23
00112e23
00912a23
01212823
01312623
0105d693
00058793
00050413
01065713
0c069c63
12071863
01061593
01079513
0105d593
01055513
8f9ea0ef
00050593
00040513
f44eb0ef
00050413
04050863
ffc52603
02400713
ffc67613
ffc60613
04c76e63
01300693
00050793
02c6f263
00052023
00052223
01b00793
06c7f463
00052423
00052623
01050793
0ce60a63
0007a023
0007a223
0007a423
01c12083
00040513
01812403
01412483
01012903
00c12983
02010113
00008067
00000593
e81eb0ef
01c12083
00040513
01812403
01412483
01012903
00c12983
02010113
00008067
00850793
0007a023
0007a223
0007a423
fa9ff06f
06071c63
00068913
00060993
01079513
01061593
0105d593
01055513
81dea0ef
00050493
01091593
01099513
0105d593
01055513
805ea0ef
0104d793
00f505b3
0105d793
02079a63
01049493
01059593
0104d493
0095e5b3
ef1ff06f
00070913
00058993
fa9ff06f
00052823
01850793
00052a23
f25ff06f
014000ef
00c00793
00f52023
00000413
f1dff06f
040017b7
9e47a503
00008067
fc010113
02c10313
02d12623
00030693
00112e23
02e12823
02f12a23
03012c23
03112e23
00612623
addfe0ef
01c12083
04010113
00008067
00050e13
04001537
fc010113
9e452503
02810313
02c12423
02d12623
00058613
00030693
000e0593
00112e23
02e12823
02f12a23
03012c23
03112e23
00612623
a8dfe0ef
01c12083
04010113
00008067
fd010113
02812423
01312e23
01612823
02112623
02912223
03212023
01412c23
01512a23
00050b13
00058993
00060413
ca4f50ef
00100793
02f51063
fff98793
0fe00713
00f76a63
0ff9f713
00e10623
00100913
02c0006f
05c40693
00098613
00c10593
000b0513
7c8040ef
fff00793
00050913
0af50463
08050e63
00c14703
00000493
fff00a13
00a00a93
0280006f
00042783
00178693
00d42023
00e78023
00148493
00c10793
009787b3
0724f463
0007c703
00842783
fff78793
00f42423
fc07d8e3
01842683
00070593
00040613
000b0513
00d7c463
fb571ce3
ca5f10ef
fd4510e3
fff00913
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00090513
02012903
03010113
00008067
00098913
fd1ff06f
00c45783
0407e793
00f41623
fc1ff06f
00c61783
01279713
02074063
06462703
000026b7
00d7e7b3
000026b7
00d76733
00f61623
06e62223
eadff06f
fe010113
040017b7
00812c23
9e47a403
00112e23
00058613
00050593
00040663
03842783
04078063
00c61783
01279713
02074063
06462703
000026b7
00d7e7b3
000026b7
00d76733
00f61623
06e62223
00040513
01812403
01c12083
02010113
e49ff06f
00a12423
00040513
00c12623
d09ea0ef
00c12603
00812583
fadff06f
ff010113
00058713
00812423
00912223
00050413
042594b7
00060593
00070513
00112623
b404a823
661040ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
01052603
4055de13
08ce5663
01450313
00261813
002e1793
01f5f593
01030833
00f307b3
06058e63
0007a683
02000e93
00478793
40be8eb3
00b6d6b3
0507f663
00030893
0007a703
00488893
00478793
01d71733
00d76733
fee8ae23
ffc7a683
00b6d6b3
ff07e0e3
41c60633
00261613
ffc60613
00c30633
00d62023
04068663
00460613
0440006f
00d52a23
00030613
fe0698e3
00052823
00052a23
00008067
00030713
ff07f8e3
0007a683
00478793
00470713
fed72e23
ff07e8e3
41c60633
00261613
00c30633
406607b3
4027d793
00f52823
fc6602e3
00008067
fa010113
00025837
05312623
92082983
05412423
03912a23
00050a13
00058c93
00098513
05212823
05512223
03812c23
03b12623
00d12423
00e12023
00f12623
04112e23
04812c23
04912a23
05612023
03712e23
03a12823
00060913
b00ec0ef
000cac03
00a986b3
03000713
002c4783
fff6cd83
00050a93
60e79e63
ffe00693
003c0813
418686b3
03000593
00084783
01068b33
00080c13
00180813
feb788e3
00025d37
820d0d13
00fd07b3
0007c783
2e078e63
000c4783
00000813
00000413
00fd07b3
0007c783
000c0493
00078c63
0014c783
00148493
00fd07b3
0007c783
fe0798e3
000a8613
00098593
00048513
01012223
2fd000ef
00412803
00050b93
12051c63
54040c63
0004c783
409406b3
00269b93
0df7f793
05000593
00048413
12b78e63
009ca023
1c081463
418407b3
fff78793
00700713
00000593
00f75863
4017d793
00158593
fef74ce3
000a0513
869f50ef
00050b13
6e050e63
01450493
00048893
568c7063
00100e93
00000c93
00000713
415e8eb3
02000e13
fff44783
fff40813
1bb78e63
21cc8663
000c8593
004c8c93
fff44783
00080413
00fd07b3
0007c803
00f87813
00b81833
01076733
fc8c66e3
00488613
40960633
40265613
00e8a023
00cb2823
00070513
00561413
b65f50ef
00092983
40a40633
26c9c863
00000c13
45364a63
00892783
4b77ca63
00492703
20ebd663
41770bb3
2b3bc663
00c92783
00200693
54d78463
00300693
52d78a63
00100693
4ed78663
000b0593
000a0513
83df50ef
00012783
05000413
0007a023
0cc0006f
0004c783
00000b93
ec040ae3
409406b3
0df7f793
05000593
00269b93
00048413
ecb796e3
00144783
02b00593
3cb78663
02d00593
1cb78863
00140893
00000313
00fd07b3
0007c583
01800513
00040493
fff58793
0ff7f793
e8f56ae3
0018c783
ff058593
00188493
00fd07b3
0007c503
01900e13
02050863
02ae4663
0014c883
00259793
00b787b3
00179793
011d05b3
00a787b3
0005c503
00148493
ff078593
fc051ce3
00030463
40b005b3
009ca023
00bb8bb3
e40800e3
01603433
40800433
ffa47413
00640413
05c12083
00040513
05812403
05412483
05012903
04c12983
04812a03
04412a83
04012b03
03c12b83
03812c03
03412c83
03012d03
02c12d83
06010113
00008067
01d807b3
e587e2e3
00078513
000a8613
00098593
01d12e23
01112c23
01012a23
00e12823
00f12223
089000ef
00412783
01012703
01412803
01812883
01c12e83
02000e13
e00512e3
00078413
de8c68e3
e25ff06f
00e8a023
00000593
00488893
00400c93
00000713
dedff06f
000a8613
00098593
000c0513
039000ef
12051c63
015c0433
00044683
00dd07b3
0007c783
12078663
03000713
00040c13
00e69c63
001c4783
001c0c13
fee78ce3
00fd07b3
0007c783
0017b813
00100b13
ccdff06f
00100413
020c0263
00c92783
00200713
10e78063
00300713
10e78463
00100713
1ee78863
01046413
00012783
0167a023
00812783
0177a023
ec9ff06f
00100313
00244783
00240893
e31ff06f
41360433
00040593
000b0513
fa4f60ef
00050c13
02050a63
fff40713
40575793
00279793
00f487b3
0007a603
00100793
00e797b3
00c7f7b3
00100c13
00078663
24ec4a63
00200c13
00040593
000b0513
a89ff0ef
008b8bb3
d45ff06f
fffb8c93
200c1863
200c9e63
405cd793
00279793
00f487b3
0007a703
00100793
019797b3
00e7f7b3
00078463
002c6c13
000b8593
000b0513
a45ff0ef
417989b3
00200413
00492b83
f15ff06f
000c4683
000c0413
0df6f693
05000793
1ef68a63
008ca023
de5ff06f
00c12703
00100793
40e787b3
00f12623
00c12783
f00780e3
010b2a83
00048793
fff00613
002a9c13
018485b3
0100006f
00478793
fe07ae23
20b7fa63
0007a703
fec708e3
00170713
00e7a023
00200793
22f40a63
01f9f993
02100413
ea098ee3
01848c33
ffcc2503
fbcf50ef
02000793
413787b3
eaf552e3
010b2783
28f05c63
014b2603
00279793
00f487b3
018b0593
00165613
26f5fa63
00048513
0005a703
00450513
00458593
01f71713
00c76733
fee52e23
ffc5a603
00165613
fef5e0e3
416787b3
fe778793
ffc7f793
00478793
00f487b3
00c7a023
24061463
40978733
40275713
00eb2823
22978863
00892783
001b8b93
0977ce63
02100413
e1dff06f
002c7793
e00788e3
0004a783
00fc67b3
0017f793
f00792e3
01046413
dfdff06f
00000313
e0dff06f
40c98433
000b0593
00040613
000a0513
cf9f50ef
00050b13
408b8bb3
01450493
b91ff06f
015485b3
0005c783
00058493
00fd0533
00054503
aa0502e3
0014c783
00148493
00fd06b3
0006c683
fe0698e3
409585b3
00259b93
a85ff06f
002c0c13
00000b13
a05ff06f
000b0593
000a0513
bb8f50ef
00012783
0a300413
0007a023
c49ff06f
00100c13
df5ff06f
00000713
aedff06f
000c8593
000b0513
d28f60ef
00050c13
dd9ff06f
ffe40593
000b0513
d14f60ef
00300c13
da0512e3
d9dff06f
00000b93
00100813
b5dff06f
b1799ce3
00f98c63
fff98593
000b0513
ce8f60ef
b00502e3
00492703
00812783
06200413
00e7a023
00100793
00fb2823
00f4a023
00012783
0167a023
bc1ff06f
00c12783
ac078ae3
fd5ff06f
00c12783
ac0794e3
fc9ff06f
008b2703
000a8793
06ead463
00478713
00271713
00178793
00eb0733
00fb2823
00100613
00c72223
00200713
00e40663
e0fac0e3
dd5ff06f
00092783
02200413
fff78793
c93794e3
4059d793
00279793
00f487b3
0007a783
00100413
01341433
00f47433
00143413
02140413
c61ff06f
004b2583
000a0513
00158593
9e0f50ef
00050c93
04050c63
010b2603
00cb0593
00c50513
00260613
00261613
f79f40ef
000b0593
000a0513
a5cf50ef
010ca783
014c8493
000c8b13
f55ff06f
00c4a023
00048793
00061863
000b2823
000b2a23
dd1ff06f
00478793
db9ff06f
000256b7
00025537
ef868693
00000613
08400593
01c50513
9f4ff0ef
000256b7
00025537
ef868693
00000613
0de00593
01c50513
9d8ff0ef
00052683
01900813
0005c603
00168693
00158593
02060263
0006c703
fbf70793
0ff7f793
00f86463
02070713
fcc70ee3
00000513
00008067
00d52023
00100513
00008067
fe010113
01212a23
0005a903
00812e23
00912c23
40595793
00279793
01312823
01412623
01f97913
00f607b3
18091863
ffc78893
00078493
00052683
fe04ae23
0016c703
1a070863
00025fb7
00088f13
00088813
00000593
00000293
00000313
820f8f93
00800413
02000393
00700993
03c0006f
16e3ec63
0262d463
01e87463
10b9d263
00800593
01067c63
ffc80f13
fe082e23
00030293
000f0813
00000593
0026c703
00168693
02070e63
00ef87b3
0007c783
fc0780e3
00158593
00130313
0ab44663
00082703
00471713
00f7f793
00e7e7b3
00f82023
0026c703
00168693
fc0716e3
10030863
01e87663
00700793
16b7d463
0d067a63
00060713
00080793
0007a683
00478793
00470713
fed72e23
fef8f8e3
00188693
00180713
00400793
12e6f463
00f607b3
00478793
fe07ae23
fef8fce3
ffc4a783
00079a63
0d160c63
ffc8a783
ffc88893
fe078ae3
01c12403
01812483
01412903
01012983
00c12a03
00500513
02010113
00008067
f3067ae3
fe082e23
00000713
ffc80813
00100593
f4dff06f
40b405b3
00082e03
00259593
40b38a33
00080793
0047ae83
00478793
014e9733
01c76733
00bede33
fee7ae23
01c7a023
ffe7e2e3
ecdff06f
00478493
00078893
e75ff06f
ffc4a783
f60906e3
02000693
412686b3
fff00713
00d75733
00e7f7b3
fef4ae23
f51ff06f
02900793
04f70663
01c12403
01812483
01412903
01012983
00c12a03
00400513
02010113
00008067
01c12403
00100793
00f8a023
01812483
01412903
01012983
00c12a03
00500513
02010113
00008067
00268693
00d52023
ea1ff06f
410887b3
ffc7f793
00478793
ed1ff06f
00800513
40b50533
00082683
00251513
02000313
40a30333
00080793
0047a583
00478793
00659733
00d76733
00a5d6b3
fee7ae23
00d7a023
ffe7e2e3
e70662e3
f31ff06f
ff010113
00812423
00912223
00050413
042594b7
00058513
00112623
b404a823
23c040ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
0ff00793
00a7ee63
000247b7
c0178793
00f50533
00054503
00857513
00008067
00000513
00008067
00000513
00008067
000257b7
1487a503
14c7a583
00008067
0a060063
00b567b3
0037f793
08079e63
00300793
08c7fa63
feff0337
808088b7
eff30313
08088893
00300e13
01c0006f
ffc60613
06060663
06079463
00450513
00458593
06ce7263
00052703
0005a683
006707b3
fff74813
0107f7b3
0117f7b3
fcd708e3
00054683
0005c803
05069a63
00050713
0140006f
00074683
0005c803
05069063
00078e63
00170713
40e607b3
fff78793
00158593
00f507b3
fc069ee3
00000513
00008067
00054683
0005c803
00d81863
00100793
faf61ce3
fe5ff06f
41068533
00008067
01052603
4055de13
08ce5663
01450313
00261813
002e1793
01f5f593
01030833
00f307b3
06058e63
0007a683
02000e93
00478793
40be8eb3
00b6d6b3
0507f663
00030893
0007a703
00488893
00478793
01d71733
00d76733
fee8ae23
ffc7a683
00b6d6b3
ff07e0e3
41c60633
00261613
ffc60613
00c30633
00d62023
04068663
00460613
0440006f
00d52a23
00030613
fe0698e3
00052823
00052a23
00008067
00030713
ff07f8e3
0007a683
00478793
00470713
fed72e23
ff07e8e3
41c60633
00261613
00c30633
406607b3
4027d793
00f52823
fc6602e3
00008067
ff010113
00812423
00058413
0105a583
01440793
00912223
00259693
00112623
01212023
00050493
00d786b3
fff00613
0100006f
00478793
fe07ae23
02d7f863
0007a703
fec708e3
00c12083
00040513
00812403
00170713
00e7a023
00412483
00012903
01010113
00008067
00842783
02f5de63
00458793
00279793
00158593
00b42823
00c12083
00f407b3
00040513
00812403
00100713
00e7a223
00412483
00012903
01010113
00008067
00442583
00048513
00158593
b6df40ef
00050913
02050a63
01042603
00c40593
00c50513
00260613
00261613
905f40ef
00040593
00048513
be9f40ef
01092583
00090413
f85ff06f
000256b7
00025537
ef868693
00000613
0c100593
07850513
ba5fe0ef
fb010113
03412c23
03812423
00070a13
00068c13
01810713
01c10693
04812423
04912223
05212023
03312e23
03512a23
03612823
03912223
05012b03
04112623
03712623
03a12023
00050913
00078a93
00080993
00088413
9f1f50ef
01812603
000c2c83
01c12303
00050493
419605b3
00658333
00b12c23
00612e23
08b05c63
03500793
02fc8a63
00100793
26f40c63
00200793
12f40463
fff58713
30071663
00000b93
02098463
01452783
0017d793
0017f793
3100006f
00000b93
00098863
00cc2703
00100793
32f70263
00090513
00048593
ae9f40ef
04c12083
04812403
04412483
04012903
03c12983
03812a03
03412a83
03012b03
02812c03
02412c83
02012d03
000b8513
02c12b83
05010113
00008067
00000b93
fa098ae3
00000d13
20059463
004c2783
06f35063
40678433
00f12e23
008cc663
010c2783
14078e63
05000793
0004a823
00fb2023
c61fe0ef
02200793
00f52023
01c12303
00000d13
006a2023
00048613
000c8593
000a8513
b81f50ef
000b2783
00100b93
01a7e7b3
00fb2023
f49ff06f
008c2783
fc67dae3
0a300713
00178793
00eb2023
00f12e23
c0dfe0ef
02200793
00f52023
01c12303
0004a823
00000d13
fa9ff06f
b9df50ef
01812583
00050b93
00048513
c49ff0ef
00048593
00090513
d19ff0ef
01fcf413
00050493
22041663
0104a783
00378793
00279793
00f487b3
0047a503
c95f40ef
22850863
000b9663
0144ab83
001bfb93
0104a603
20c05a63
0144a683
01448593
00261613
00c58633
01848793
0016d693
1ec7f663
0007a703
00478793
01f71713
00d76733
ffc7a683
fee7ac23
0016d693
fec7e2e3
409607b3
fe778793
ffc7f793
00478793
00f587b3
00d7a023
1c069863
40b78733
40275713
00e4a823
00f59463
0004aa23
01c12303
02000d13
00130313
00612e23
e91ff06f
fff40c13
0a0c0c63
0a0b8263
405c5793
00478793
00279793
00f487b3
0047a703
00100793
018797b3
00040593
00048513
00e7f433
b49ff0ef
00200793
00fb2023
05000d13
0a040c63
00048593
00090513
c09ff0ef
00050493
abdfe0ef
02200793
00f52023
06000d13
0940006f
a55f50ef
01812583
00050b93
00048513
b01ff0ef
01703433
01c12303
00441d13
e01ff06f
00050593
40cc8633
00090513
968f50ef
01c12303
00050493
de5ff06f
000c0593
00048513
a0df50ef
00050b93
f40b98e3
d6098ae3
405c5793
00478793
00279793
00f487b3
0047a703
00100793
018797b3
00040593
00048513
00e7f433
a91ff0ef
00200793
00fb2023
f40418e3
a19fe0ef
02200793
00f52023
01c12303
dbdff06f
40575793
00478793
00279793
00f507b3
0047a783
00e7d7b3
0017f793
00048513
00f12623
98df50ef
01812583
00050b93
00048513
a39ff0ef
00c12783
f2078ae3
de9ff06f
96df50ef
01812583
00a03433
00050b93
00048513
a15ff0ef
01c12303
00441d13
d19ff06f
02000793
40878433
dd1ff06f
00d4aa23
00058793
00069c63
0004a823
e55ff06f
01c12303
02000d13
cedff06f
00478793
e31ff06f
01052703
01450513
fff00693
00271713
00e50733
0100006f
00450513
fed52e23
00e57a63
00052783
fe0788e3
fff78793
00f52023
01000513
00008067
ff010113
0045a783
00912223
01f60493
00812423
00112623
01212023
4054d493
00060413
00058693
0a97c263
01f47513
01468593
40545413
06051e63
00241713
0086a823
00e58733
04e5f863
00058793
fff00613
00478793
fec7ae23
fee7ece3
01568793
00400613
00f76a63
40d707b3
feb78793
ffc7f793
00478613
00c585b3
00050c63
ffc5a783
02000713
40a70733
00e7d7b3
fef5ae23
00c12083
00812403
00412483
00012903
00068513
01010113
00008067
00140413
00241713
0086a823
00e58733
f8e5e4e3
fbdff06f
00050913
e6cf40ef
00048593
00090513
db8f40ef
00050693
f40514e3
000256b7
00025537
ef868693
00000613
10000593
07850513
e20fe0ef
f2010113
000258b7
0d612023
9208ab03
0c812c23
0d212823
00050413
00068913
000b0513
0c912a23
0d412423
0b812c23
00058a13
0ba12823
02d12423
04e12823
02f12c23
0c112e23
0d312623
0d512223
0b712e23
0b912a23
0bb12623
00c12c23
00080493
ed1ea0ef
00092c03
000257b7
00050d13
08012423
08012c23
000a0713
02d00593
92c78693
08e12a23
00074783
00070913
00f5ea63
00279613
00d60633
00062603
00060067
04012023
03000713
00000c93
1ee78a63
02812683
02f00713
00078d93
0106a683
06d12223
1ef778e3
00090513
00000a93
00000993
00000493
03900693
00800593
00f00813
02f00613
13b6c263
1095c263
00299713
013709b3
00199993
00f989b3
fd098993
00150513
08a12a23
00054d83
00148493
000d8793
fdb648e3
000d0613
000b0593
e9cff0ef
00048b93
1a0518e3
09412783
00012e23
01a787b3
08f12a23
0007cd83
fd0d8613
00900793
16c7e0e3
09412803
00150513
00060d93
00060463
7cc0106f
00180793
08f12a23
00184d83
fd5ff06f
00100793
04f12023
00170913
09212a23
00174783
f0079ee3
00600793
08f12423
01812783
00600513
00078863
01812783
0147a023
08812503
0dc12083
0d812403
0d412483
0d012903
0cc12983
0c812a03
0c412a83
0c012b03
0bc12b83
0b812c03
0b412c83
0b012d03
0ac12d83
0e010113
00008067
00170713
e95ff06f
f0984ae3
002a9713
01570ab3
001a9a93
00fa8ab3
fd0a8a93
efdff06f
000d0613
000b0593
dacff0ef
0c051263
09412783
01a787b3
08f12a23
0007cd83
00048463
1950106f
03000713
00ed8463
0610106f
00100713
40f70733
03000693
00e78533
00178793
08f12a23
0007cd83
fedd88e3
fcfd8793
00800713
02f76ce3
09412903
00150793
fd0d8d93
00f12e23
00090813
00000b93
00100493
00299793
013787b3
00179793
00fd89b3
00000513
ec9ff06f
00194783
05800613
00190713
0df7f793
03000693
00c79463
5340106f
08e12a23
00074783
00070913
00170713
fed788e3
0e078e63
00100c93
dd9ff06f
00048b93
00000513
00012e23
00000713
fdfdf793
04500693
00000b13
08d79463
00a4e7b3
0197e7b3
0a078e63
09412a03
02b00793
001a0693
08d12a23
001a4d83
00fd9463
4740106f
02d00793
00000693
00fd9a63
00100693
002a0793
08f12a23
002a4d83
fd0d8793
00900613
7af66463
03000793
02fd9063
09412783
03000613
00178793
08f12a23
0007cd83
00178793
fecd8ae3
fcfd8793
00800613
00000b13
20f670e3
0a049263
00ace533
04051263
02071a63
06900793
28fd82e3
09b7c063
04900793
26fd8ce3
04e00793
00fd9c63
000255b7
fd858593
09410513
888ff0ef
2a051ee3
00600793
08f12423
09412a23
01812703
00070663
09412783
00f72023
04012783
09812603
00078863
08812783
0087e793
08f12423
da060ae3
03812503
000c0593
b64f50ef
09812583
00040513
a24f40ef
08812503
d99ff06f
06e00793
f8fd88e3
fa1ff06f
02812783
01c12683
00100713
00c7a783
40db06b3
04d12423
04012683
0037f793
08e12423
40d78633
00200713
02c12a23
00e78e63
00168693
00300713
02d12a23
00e78663
0017b793
02f12a23
000b9463
00048b93
01000793
00048a13
0097d463
01000a13
00098513
388060ef
00900793
00050313
00058e13
0497d863
ff7a0793
00024737
f6870713
00379793
00e787b3
0007a603
0047a683
2ac050ef
00050c93
000a8513
00058a93
348060ef
00050613
00058693
000c8513
000a8593
078040ef
00050313
00058e13
03500c93
0d8cce63
00f00793
0c97ca63
04812703
00071463
5bc0106f
04812683
00d04463
5fc0106f
01600713
00d74463
6ec0106f
04812683
02500713
41448cb3
40970733
00dc8cb3
0ad74463
40978ab3
00024cb7
f68c8c93
003a9793
019787b3
0007a503
0047a583
00030613
000e0693
20c050ef
04812783
415787b3
00379793
019787b3
0007a603
0047a683
1f0050ef
08810793
00f12023
03412883
03812783
05012703
02812683
00050313
00058e13
00058613
00000813
00050593
00040513
02612023
01c12a23
cc0ff0ef
01412e03
02012303
e00516e3
00000c93
0080006f
04812c83
41448a33
019a0cb3
53905263
00fcf793
02078863
00024737
f6870713
00379793
00e787b3
0007a503
0047a583
00030613
000e0693
164050ef
00050313
00058e13
ff0cfc93
620c9c63
00030893
000e0813
08c10713
00088593
09010693
00080613
00040513
e89f40ef
09012783
08c12703
08a12c23
00fc8cb3
09912823
418705b3
00050a13
00b05c63
00bc8cb3
a2cff0ef
000c0713
09812623
09912823
02812603
00ec86b3
418686b3
00862783
04d12c23
00178793
00d7d463
7e40106f
00462783
02f12e23
00f6c463
2780106f
40fc8ab3
75504a63
020a8863
00ea8ab3
09512623
01505463
52c0106f
fff00793
00fad463
3b00106f
00100793
08f12623
00fa2823
00fa2a23
03c12703
06412783
08e12823
00079463
2340106f
05812783
00100693
00d12a23
00178793
04e12c23
00e7d463
36c0106f
00048693
00098713
000b8613
00090593
00040513
8b4f40ef
00025737
0d872683
0dc72703
04812603
06d12823
06e12a23
00025737
10072683
10472703
fff64793
06d12423
06e12623
00025737
10872683
10c72703
41f7d793
06d12c23
01c12683
06e12e23
41f65713
41668b33
00eb7733
00f677b3
00050d13
02e12023
04f12623
00000493
01812e23
004d2583
00040513
df5f30ef
00050c93
00051463
6780106f
010d2603
00cd0593
00c50513
00260613
00261613
b89f30ef
09812783
00040513
0047a583
dc1f30ef
00050913
00051463
6280106f
09812583
00c50513
0105a603
00c58593
00260613
00261613
b51f30ef
09012c03
08c12a83
00100593
00040513
a58f40ef
009c0a33
409a8bb3
00050993
180a4ae3
02012783
01478b33
04c12a03
01c12703
018a8ab3
00170793
40ea8ab3
03c12703
417787b3
00ead663
40ea8ab3
015787b3
00fb0ab3
00fa0a33
000a8793
015a5463
000a0793
00fb5463
000b0793
00f05863
40fa8ab3
40fa0a33
40fb0b33
02012783
02f05e63
00078613
00098593
00040513
d30f40ef
00090613
00050593
00050993
00040513
a70f40ef
00050c13
00090593
00040513
d85f30ef
000c0913
409a8633
0cc04ee3
460610e3
04812783
48f04e63
49404063
01605c63
00098593
000b0613
00040513
e34f40ef
00050993
000c8613
00090593
00040513
809f40ef
01052703
00100793
00050a13
00e7c863
01452783
00079463
7fd0006f
00ca2483
00098593
000a2623
000a0513
f80f40ef
03412783
5a078e63
22a052e3
00098593
000a0513
ce1f40ef
06812603
06c12683
00050b13
00058a93
539040ef
06a044e3
24048ce3
07012783
07412703
04012223
00078b13
02f12223
02000793
00070b93
02e12623
04f12a23
00000493
00000c13
08c12603
09012783
00f607b3
02f12823
01412783
00079663
01c12783
3af648e3
000b8613
08410713
08010693
000b0593
00040513
b05f40ef
08012603
00050d93
2c0644e3
340610e3
09812a83
010aa783
640c0c63
00378793
00279793
00fa87b3
0047a503
f1df30ef
09812583
000d8613
00040513
f00f40ef
01412703
08a12c23
010aa783
02071663
01052683
fff78713
48d74ee3
05812783
03c12703
08e79ce3
08c12783
01812a23
fff78793
08f12623
000d8593
00040513
bf5f30ef
000a8593
00040513
be9f30ef
6a049ee3
08c12703
09012783
00e787b3
03012703
18e78ce3
01412783
08078ce3
00090593
00040513
bbdf30ef
000c8593
00040513
bb1f30ef
00098593
00040513
ba5f30ef
000a0593
00040513
b99f30ef
cf1ff06f
00000b93
00012e23
00000493
00100713
83dff06f
000d0613
000b0593
00090513
d01fe0ef
00051463
7dd0006f
00000b93
00000a93
00000993
00000493
00000513
00012e23
00000713
00000b13
895ff06f
09412a23
00000b13
889ff06f
b00c8ee3
41900cb3
00fcf793
02078863
00024737
f6870713
00379793
00e787b3
0007a603
0047a683
00030513
000e0593
208040ef
00050313
00058e13
ff0cfc93
ac0c8ee3
404cdd93
00f00713
01b74463
2880106f
00024737
801007b7
05072a03
05472a83
fff78793
00000693
00f12a23
000d8c93
00068793
00030513
01412703
3ff006b7
c0178793
00ee7733
00d76733
014e5e13
7ffe7e13
00050613
00070693
000a0513
000a8593
00fe0d33
3c1040ef
ff0c8c93
00f00713
000d0793
00058e13
fb974ee3
00050313
00fdfd93
014e5c93
801006b7
7ffcfc93
fff68693
00de76b3
c01c8c93
3ff00e37
01ac8cb3
01c6ee33
a20d86e3
00024d37
00030a93
000e0a13
030d0d13
00030893
00000693
000e0593
001df793
00078e63
004d2683
000d2603
00088513
349040ef
00050893
00100693
401ddd93
008d0d13
fc0d9ce3
00058813
9e0692e3
000a8893
000a0813
9d9ff06f
404cdd93
00f00793
01b7c463
7a90006f
000247b7
0787aa03
07c7aa83
801007b7
fff78793
00000693
00f12a23
000d8c93
00068793
00030513
01412703
3ff006b7
c0178793
00ee7733
00d76733
014e5e13
7ffe7e13
00050613
00070693
000a0513
000a8593
00fe0d33
2b5040ef
ff0c8c93
00f00713
000d0793
00058e13
fb974ee3
00050313
00fdfd93
014e5c93
801006b7
7ffcfc93
fff68693
00de76b3
c01c8c93
3ff00e37
01ac8cb3
01c6ee33
920d80e3
00024d37
00030a93
000e0a13
058d0d13
00030893
00000693
000e0593
001df793
00078e63
004d2683
000d2603
00088513
23d040ef
00050893
00100693
401ddd93
008d0d13
fc0d9ce3
ef5ff06f
000c8593
000a0613
00040513
9bcf40ef
00050c93
b71ff06f
04c12603
000c8593
00040513
84cf40ef
00050c93
b5405ce3
fd1ff06f
09412803
fd0d8b13
02f00893
00180793
08f12a23
00184d83
03900613
02f00593
13b8da63
03b64663
002b1893
016888b3
00078313
00178793
00189893
08f12a23
01b888b3
00134d83
fd088b13
fdb5cce3
410787b3
00800613
0ef65e63
00005b37
e1fb0b13
da068063
41600b33
d98ff06f
04012023
b8cff06f
000a8613
000a0593
00040513
910f40ef
08c12783
08a12c23
015787b3
08f12623
8c1ff06f
000255b7
fcc58593
09410513
e1cfe0ef
d8050c63
09412783
000255b7
fd058593
fff78793
09410513
08f12a23
dfcfe0ef
00051863
09412783
00178793
08f12a23
02812783
00300713
08e12423
0087a783
05012703
00178793
00f72023
d58ff06f
02812783
05012703
0087a783
00178793
00f72023
09412783
0007c703
00400793
08f12423
02800793
d2f71663
02812483
03812603
09410513
00048593
dd0fe0ef
0084a783
05012703
08a12423
00178793
00f72023
d00ff06f
000057b7
e1f78793
f167d4e3
00078b13
f01ff06f
2e054ee3
a40514e3
01c12c03
460480e3
01412783
140782e3
08c12603
09812583
fff00513
40565693
01458793
00269693
00d786b3
66d7f4e3
0007a703
00478793
fea70ae3
01100793
08f12423
5b8bdce3
0145a783
0017f793
04078a63
00040513
a21fe0ef
01052703
08c12483
08a12c23
00370713
00271713
00e507b3
0047a503
409004b3
01f4f493
999f30ef
00950863
08c12783
00178793
08f12623
02100793
08f12423
01412783
0c0788e3
09012783
05012703
00090593
00040513
00f72023
e8cf30ef
000c8593
00040513
e80f30ef
00098593
00040513
e74f30ef
000d0593
00040513
e68f30ef
000a0593
00040513
e5cf30ef
02812783
09012703
0087a783
3ce7cce3
06412703
09812783
58071863
0107a783
08812703
00f027b3
ff877713
00179793
03077693
00e7e7b3
00068463
0407e793
08f12423
805fd0ef
02200793
00f52023
ba4ff06f
010da703
46e7d463
000a8e13
000d8793
0047a583
00040513
07c12023
04f12e23
d3cf30ef
05c12783
06012e03
00050c13
5e050ae3
0107a383
01450893
00010eb7
007c2823
010e2603
01478513
014e0e13
00261593
00b885b3
00050f13
00088313
00000793
fffe8e93
000f2703
000e2803
00430313
01d776b3
01d87fb3
01f686b3
00f686b3
01085813
01075793
010787b3
0106d713
00e787b3
01079713
01d6f6b3
00d76733
fee32e23
004f0f13
004e0e13
0107d793
fab36ae3
015c0693
00400713
00d5ea63
41858733
feb70713
ffc77713
00470713
40c38633
00261613
00c58633
00e888b3
00e505b3
04c8f263
00010537
fff50513
0005a683
00488893
00458593
00a6f733
00f70733
01075793
0106d693
00d787b3
01079693
00a77733
00e6e733
fee8ae23
0107d793
fcc8e6e3
34079663
010aa783
fff38393
09812c23
36f3c663
01412783
46078463
08c12783
01c12703
00178793
40e78733
08f12623
00e037b3
00f12a23
8a5ff06f
00090593
00040513
d75f30ef
00050913
f1cff06f
04c12783
02012b03
41478a33
e70ff06f
000257b7
0f87a603
0fc7a683
000b0513
000a8593
59c040ef
02a12223
02b12623
34048a63
01000793
04f12a23
00000c13
02412a83
02c12483
07812603
07c12683
000a8513
00048593
484040ef
32055c63
00048593
000a8513
460050ef
04a12223
554050ef
00058b93
00050613
00050b13
00048593
000a8513
000b8693
401040ef
03412703
00100793
02a12223
02b12623
02f70463
00200793
4ef70463
000257b7
0f87a603
0fc7a683
340040ef
02055063
00000493
f18ff06f
fe0c0ce3
00000613
00000693
324040ef
fea054e3
04412783
05412703
00000493
00178793
04f12223
00078513
03000793
40e787b3
04f12a23
4c4050ef
00050b13
00058b93
ed0ff06f
09812583
00100613
00040513
c4df30ef
09012783
00050713
000d8593
fff78793
00040513
08f12823
08e12c23
b4cf30ef
05812783
000a8593
00040513
fff78793
04f12c23
b34f30ef
09812783
00000493
0107a683
01478793
00269693
00d786b3
00d7ea63
02c0006f
00478793
02048493
02d7f063
0007a703
fe0708e3
00d7fa63
09c10513
08e12e23
e3cf30ef
00a484b3
00012a23
f20ff06f
0017f793
0097cc33
16978ce3
38049863
01100793
08f12423
03c12703
05812783
02e78c63
01c12a83
01f00793
09812583
4157de63
01458793
01f00693
0140006f
fe0a8a93
00148493
00478793
4156d263
0007a703
fe0706e3
000c0493
01412783
1e078663
00100793
1777d8e3
09012703
08c12783
07012683
01412c03
00f707b3
02f12823
07412783
00068b13
04012223
00078b93
02f12623
01000793
02d12223
04f12a23
db0ff06f
04412783
e6078463
000257b7
1507a603
1547a683
000b0513
000b8593
354040ef
000257b7
02c12a83
0f87a603
0fc7a683
00050b93
02412503
00058b13
000a8593
1fd040ef
800007b7
0167c7b3
000b8613
00078693
00050d93
00058c13
230040ef
20055a63
02412603
000b8513
000a8693
000b0593
218040ef
de055a63
08812783
05412703
01c12c03
00e7e7b3
08f12423
b01ff06f
40c005b3
bf8fe0ef
d38ff06f
000d8e13
000a8793
b9dff06f
008c2783
28f38e63
00438793
00138713
00279793
00ec2823
00fc07b3
00100713
00e7a223
010aa783
09812c23
c8f3dee3
00438393
00239393
007c0c33
004c2503
04712e23
c1cf30ef
05c12383
00050c13
007a83b3
0043a503
c08f30ef
c6ac46e3
d30ff06f
00050593
00040513
a01f30ef
00050d93
cb4ff06f
415485b3
00090513
b64fe0ef
b98ff06f
02000793
04f12a23
00100c13
cb1ff06f
02412b03
02c12b83
04012223
00000493
c38ff06f
09812583
40c78db3
000d8613
00040513
00078a93
9adf30ef
09012783
08a12c23
09512623
41b787b3
08f12823
c28ff06f
0007a823
05000793
08f12423
a94fd0ef
02200793
00f52023
e35fe06f
08c12603
09012783
07012703
04012223
00f607b3
02f12823
07412783
00070b13
02e12223
00078b93
02f12623
01000793
04f12a23
00100c13
bc8ff06f
09812583
0105a703
14e05663
0145a783
01458513
00271713
00e50633
01858693
0017d793
12c6f263
0006a703
00468693
01f71713
00f767b3
fef6ac23
ffc6a783
0017d793
fec6e2e3
40b60733
fe770713
ffc77713
00470713
00e50733
00f72023
3a079063
40a707b3
4027d793
00f5a823
0ee50463
05812783
04012223
00178793
04f12c23
09012783
00178793
08f12823
bccff06f
000b8613
000d8513
000b0693
000c0593
725030ef
bea05263
000257b7
0d87a503
0dc7a583
000b8613
000b0693
79c040ef
02412603
02c12683
6fd030ef
baa05e63
dc9ff06f
00378793
00279793
00f50533
00452503
04f12e23
a40f30ef
05c12783
00050713
04e12e23
00fa87b3
0047a503
a28f30ef
05c12703
b2e54a63
b4cff06f
000257b7
0d87ab03
0dc7ab83
02100793
08f12423
02000793
000c0493
04012223
03612223
03712623
04f12a23
00000c13
a68ff06f
00f5aa23
00050713
2a079863
0005a823
0005aa23
f19ff06f
b20c0ee3
00000493
a44ff06f
004c2583
00040513
00158593
e39f20ef
00050793
6c050e63
010c2603
00cc0593
00c50513
00260613
00261613
04f12e23
bcdf20ef
000c0593
00040513
eb1f20ef
05c12783
0107a383
00078c13
d1dff06f
00000693
b9dfe06f
01c12a83
00100793
6357dc63
01458593
00249513
00a58533
9c8f30ef
fffa8a93
bf5546e3
01c12c03
09812583
05812783
000c0613
fff78793
00040513
08f12823
09812623
f14fe0ef
08a12c23
fa0ff06f
04012783
05012683
02812603
00048813
09810713
09410593
00040513
bc8fd0ef
08a12423
00600793
00f50463
bb5fe06f
01812783
09412a23
09812603
00079463
bc9fe06f
01812783
0147a023
bbdfe06f
01100793
08f12423
018bcc63
09812583
0145a703
00058793
00177713
4a071063
08c12783
00f12a23
01412783
40fc04b3
14fc1063
09012783
05012703
00090593
00040513
00f72023
dadf20ef
000c8593
00040513
da1f20ef
00098593
00040513
d95f20ef
000d0593
00040513
d89f20ef
000a0593
00040513
d7df20ef
02812783
00000493
0087a703
09012783
00f74463
b01fe06f
0a300793
08f12423
09812783
0007a823
f41fc0ef
02200793
00f52023
02812783
05012703
0087a783
00178793
00f72023
ee049463
ac9fe06f
01c12c03
e7cff06f
00012a23
df1fe06f
03c12783
04f12c23
00100793
00f12a23
dddfe06f
01c12583
00148793
00100693
00a585b3
00b12e23
00078713
04d50c63
009505b3
00048713
00800513
fff58593
01000893
00078493
02e56263
00299693
013689b3
00199993
02f58463
00178793
00048713
00078493
fee572e3
fef8c6e3
002a9693
01568ab3
001a9a93
fddff06f
00270713
00800793
0a97c463
00070493
8e1fe06f
09812503
22905063
00050593
00048613
00040513
d50f30ef
08a12c23
09012783
409787b3
08f12823
ea1ff06f
00470713
c61ff06f
01c12c03
1c049663
02100793
08f12423
00100793
d977ca63
01412783
d8079a63
05812783
03c12703
e4e78ae3
000a0593
00100613
00040513
cf8f30ef
00098593
00050a13
e7cf30ef
e2a05ae3
09812583
01100793
08f12423
09012783
000c0613
418787b3
d91ff06f
01000793
1ae7c463
002a9793
015787b3
00179793
00f60ab3
00070493
00000513
efcfe06f
09812a03
05012783
03c12703
000a2823
000a2a23
00e7a023
05000793
08f12423
d95fc0ef
02200793
00f52023
d50ff06f
00000513
fc0fe06f
09412783
00000993
00000a93
01a787b3
08f12a23
0007cd83
f78fe06f
08810793
00f12023
03412883
03812783
05012703
02812683
000e0613
00030593
00100813
00040513
02612023
01c12a23
f85fd0ef
01412e03
02012303
00050463
8cdfe06f
00000c93
ac9fe06f
04812703
fea00793
00070c93
00f75463
ab5fe06f
01c12783
00024737
f6870713
416787b3
00379793
00e787b3
0007a603
0047a683
00030513
000e0593
1ec030ef
a31fe06f
00100793
1efb8a63
02100793
08f12423
1d8bda63
01412783
ce078ae3
09812783
0147a703
00177713
c0070c63
0107a683
01478793
fff00613
00269693
00d786b3
0100006f
00478793
fec7ae23
00d7fa63
0007a703
fe0708e3
fff70713
00e7a023
01100793
08f12423
bd0ff06f
00100493
d11ff06f
00048b93
00012e23
d78fe06f
01412783
418785b3
cb1fd0ef
dedff06f
03c12783
000a0513
419785b3
c9dfd0ef
ae5fe06f
00070493
00000513
d68fe06f
00000d13
8d0ff06f
000257b7
00269713
9e478793
00e787b3
08612e23
0007aa83
18031a63
001007b7
00fe67b3
09c10513
02612023
01c12a23
08f12e23
d41f20ef
02012303
01412e03
01500c93
40ac8cb3
04812783
00024737
f6870713
00379793
00e787b3
0007a503
0047a583
00030613
000e0693
2f5030ef
08810793
00f12023
03412883
03812783
05012703
02812683
019a8833
00050313
00058e13
00058613
03682813
00050593
00040513
02612023
01c12a23
dc1fd0ef
00050463
f10fe06f
01412e03
02012303
00000c93
905fe06f
40f007b3
ff07f793
02178793
01c12c03
08f12423
aa4ff06f
0145a703
00058793
00177713
a8070e63
a4049463
00100713
e6eb9ee3
03c12783
0005a823
08f12823
05000793
08f12423
b09fc0ef
02200793
00f52023
a64ff06f
01c12c03
09812583
fd5ff06f
09812783
0147a703
00177713
a4070463
e39ff06f
05812783
03c12703
09712423
09812583
cee790e3
0105a783
02100713
08e12423
a3779063
0145a783
a1779c63
00100793
06f12223
a0cff06f
01f67713
06071063
03c12783
00100713
00e5a823
00fc07b3
fff78793
08f12823
02100793
00e5aa23
08e12623
08f12423
ab5ff06f
09c10513
03c12023
00612a23
bbdf20ef
01412303
02012e03
40ac8cb3
e81ff06f
00000d13
df1fe06f
01c12c03
9e9ff06f
0007a603
fff00693
00e697b3
00c7e7b3
f8d78ae3
930ff06f
000256b7
00025537
ef868693
00000613
31d00593
07850513
801fc0ef
000256b7
00025537
ef868693
00000613
31b00593
07850513
fe4fc0ef
000256b7
00025537
ef868693
00000613
06a00593
07850513
fc8fc0ef
000256b7
00025537
ef868693
00000613
04200593
07850513
facfc0ef
0a300793
000a2823
08f12423
9a9fc0ef
02200793
00f52023
02812783
05012703
0087a783
00178793
00f72023
d34fe06f
00862783
fd010113
01312e23
01412c23
02112623
02812423
02912223
03212023
01512a23
01612823
01712623
01812423
00062983
00060a13
14078863
0085a783
0005a703
00050a93
00058493
0d40006f
00c4d783
4807f693
08068a63
0144a603
0104a583
00161693
00c686b3
40b70433
01f6db13
00db0b33
00140713
401b5b13
01270733
000b0613
00eb7663
00070b13
00070613
4007f793
0a078a63
00060593
000a8513
ee5e70ef
00050c13
0a050e63
0104a583
00040613
becf20ef
00c4d783
b7f7f793
0807e793
00f49623
408b0733
008c0533
0164aa23
0184a823
00a4a023
00090b13
00e4a423
00090413
00040613
000b8593
cd8f20ef
0084a783
0004a703
008a2683
416787b3
00870733
00f4a423
00e4a023
412686b3
00da2423
06068663
0049a903
0009ab83
00078b13
00898993
00078413
00070513
fe0904e3
f0f97ae3
00090b13
00090413
fa5ff06f
000a8513
8c9f30ef
00050c13
f6051ae3
0104a583
000a8513
90de70ef
00c4d783
00c00713
00eaa023
0407e793
00f49623
000a2423
fff00513
0080006f
00000513
02c12083
02812403
000a2223
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
00c5d783
ed010113
11412c23
11612823
0fb12e23
12112623
12812423
12912223
13212023
11312e23
11512a23
11712623
11812423
11912223
11a12023
0807f793
00d12423
00058a13
00050b13
00060d93
00078663
0105a783
680784e3
00025737
04c10a93
00000813
a4070713
00025c37
000254b7
000d8913
05512023
04012423
04012223
00012823
00012c23
00012e23
02012023
00012223
00e12623
bacc0c13
bbc48493
00080993
000a8d93
00094703
1e070e63
00090413
02500693
2ad70863
00144703
00140413
fe071ae3
41240bb3
1d240e63
04412703
017989b3
012da023
00170713
017da223
05312423
04e12223
00700693
008d8d93
28e6c263
00412783
00044703
017787b3
00f12223
1a070063
00000693
00144603
00140913
02010da3
fff00e93
00012023
05a00b93
00900c93
02a00d13
00068413
00190913
fe060793
04fbe863
00c12703
00279793
00e787b3
0007a783
00078067
00012023
fd060793
00012683
00094603
00190913
00269713
00d70733
00171713
00e787b3
00f12023
fd060793
fcfcfee3
fe060793
fafbfce3
00040693
10060c63
08c10623
02010da3
00100b93
00100c93
08c10413
00000e93
0026ff93
000f8463
002b8b93
0846ff13
04412703
000f1863
00012783
41778d33
05a04ee3
03b14603
02060863
03b10613
00cda023
00170713
00100613
00198993
00cda223
05312423
04e12223
00700613
008d8d93
18e64c63
020f8863
03c10613
00cda023
00170713
00200613
00298993
00cda223
05312423
04e12223
00700613
008d8d93
12e64ee3
08000613
5acf0a63
419e8d33
6ba04c63
019989b3
00170713
008da023
019da223
05312423
04e12223
00700613
008d8793
76e64c63
0046f693
00068863
00012703
41770cb3
139048e3
00012403
01745463
000b8413
00412783
008787b3
00f12223
76099863
00094703
04012223
000a8d93
e00716e3
50099ce3
00ca5783
0407f793
580796e3
12c12083
12812403
00412503
12412483
12012903
11c12983
11812a03
11412a83
11012b03
10c12b83
10812c03
10412c83
10012d03
0fc12d83
13010113
00008067
000b0513
01d12a23
995f10ef
00452783
00078513
02f12023
bbde80ef
00050793
000b0513
00f12e23
975f10ef
00852703
01c12783
01412e83
00e12c23
28079ee3
00094603
df9ff06f
00094603
02046413
dedff06f
00012703
00f12423
40e00733
00e12023
00094603
00446413
dd1ff06f
41240bb3
d72412e3
00044703
d95ff06f
04010613
000a0593
000b0513
ab9ff0ef
f20512e3
04812983
000a8d93
d65ff06f
04010613
000a0593
000b0513
03d12623
02d12423
03e12223
01f12a23
a89ff0ef
ee051ae3
04812983
04412703
02c12e83
02812683
02412f03
01412f83
000a8d93
e2dff06f
00812783
00040693
02010da3
0007a403
00478d13
3a0400e3
fff00713
00d12a23
2cee82e3
000e8613
00000593
00040513
01d12423
e09f10ef
00812e83
01412683
400506e3
40850cb3
01a12423
00000e93
0980006f
00812783
00040693
02010da3
0007a703
00478793
00f12423
08e10623
00100b93
00100c93
08c10413
d51ff06f
00040693
0206f713
1c070a63
00812783
00778793
ff87f793
0047a603
0007ac83
00878793
00f12423
00060b93
1e064263
fff00613
00068d13
00ce8863
017ce633
f7f6fd13
7a060a63
060b98e3
00900693
0796e4e3
030c8713
0ee107a3
000d0693
00100c93
0ef10413
000e8b93
019ed463
000c8b93
03b14703
00e03733
00eb8bb3
cd1ff06f
00812783
ffff86b7
8306c693
0007ac83
02d11e23
00478793
000256b7
00f12423
ea468793
00000b93
00246d13
00f12823
00200613
00000693
02d10da3
fff00693
16de8a63
017ce5b3
f7fd7693
4e059a63
260e9263
72061463
001d7c93
0f010413
f80c82e3
03000713
0ee107a3
0ef10413
f75ff06f
00812783
02047713
00478613
080716e3
01047713
200718e3
04047713
260712e3
20047693
200680e3
00812783
00c12423
0007a703
00412783
00f70023
b19ff06f
00094603
08046413
b99ff06f
00094603
06c00793
1af608e3
01046413
b85ff06f
00094603
06800793
1af606e3
04046413
b71ff06f
01046d13
020d7713
6a070a63
00812783
00100613
00778793
ff87f793
0007ac83
0047ab83
00878793
00f12423
f21ff06f
01046693
0206f713
6c070863
00812783
00778793
ff87f793
0007ac83
0047ab83
00878793
00f12423
bff6fd13
00000613
eedff06f
01046693
0206f713
e2071ae3
00812783
0106f613
0007a703
00478793
00f12423
62061463
0406f613
60060c63
01071c93
410cdc93
41fcdb93
000b8613
e20652e3
00068d13
02d00693
01903633
417008b3
02d10da3
fff00693
40c88bb3
41900cb3
00100613
e8de9ae3
00100693
e0d606e3
00200693
10d60463
0f010413
01db9793
007cf693
003cdc93
03068693
0197ecb3
003bdb93
fed40fa3
017ce7b3
00040593
fff40413
fc079ce3
001d7713
10070263
03000713
0ee68e63
ffe58593
0f010793
fee40fa3
40b78cb3
000d0693
00058413
dc9ff06f
00094603
00190713
15a602e3
fd060793
00070913
00000e93
a2fce0e3
00094603
002e9713
01d70eb3
001e9e93
00fe8eb3
fd060793
00190913
fefcf2e3
9fdff06f
02b00793
00094603
02f10da3
9e9ff06f
00812783
0007a703
00478793
00e12023
be0746e3
00094603
00f12423
9c9ff06f
00094603
00146413
9bdff06f
03b14783
00094603
9a0798e3
02000793
02f10da3
9a5ff06f
00100593
0ab600e3
00200593
00068d13
f0b610e3
01012683
0f010413
00fcf793
00f687b3
0007c703
004cdc93
01cb9793
0197ecb3
004bdb93
fee40fa3
017ce7b3
fff40413
fc079ce3
0f010793
40878cb3
000d0693
cddff06f
00012783
41778d33
a5a054e3
01000613
0ba65063
00812a23
00098793
000a0413
01000893
000d0a13
00700f13
00090d13
000e8993
00068913
00c0006f
ff0a0a13
0548da63
01078793
00170713
009da023
011da223
04f12423
04e12223
008d8d93
fcef5ee3
04010613
00040593
000b0513
de0ff0ef
3e051663
01000893
ff0a0a13
04812783
04412703
000a8d93
00700f13
fb48cae3
00090693
000d0913
000a0d13
00040a13
01412403
00098e93
00078993
01a989b3
00170713
009da023
01ada223
05312423
04e12223
00700613
008d8d93
98e650e3
04010613
000a0593
000b0513
03d12223
00d12a23
d68ff0ef
9c051ae3
02412e83
04812983
04412703
419e8d33
01412683
000a8d93
95a058e3
01000613
09a65863
00812a23
01000893
000a0413
00700e93
000d0a13
00090d13
00068913
00c0006f
ff0a0a13
0548da63
01098993
00170713
009da023
011da223
05312423
04e12223
008d8d93
fceedee3
04010613
00040593
000b0513
ce8ff0ef
2e051a63
01000893
ff0a0a13
04812983
04412703
000a8d93
00700e93
fb48cae3
00090693
000d0913
000a0d13
00040a13
01412403
01a989b3
00170713
009da023
01ada223
05312423
04e12223
00700613
008d8d93
88e65ce3
04010613
000a0593
000b0513
00d12a23
c7cff0ef
8e0514e3
04812983
04412703
01412683
000a8d93
86dff06f
04010613
000a0593
000b0513
00d12a23
c50ff0ef
8a051ee3
04812983
01412683
000a8793
869ff06f
04010613
000a0593
000b0513
c2cff0ef
88051ce3
04812983
87dff06f
00068d13
c71ff06f
01000613
0da65c63
000d0593
00090613
000d8793
000b8d13
000c8d93
00068b93
000a0913
00098693
01000893
00040993
00700293
01f12a23
03e12223
000e8c93
00060a13
00058413
00c0006f
ff040413
0488da63
01068693
00170713
0187a023
0117a223
04d12423
04e12223
00878793
fce2dee3
04010613
00090593
000b0513
b94ff0ef
4a051263
01000893
ff040413
04812683
04412703
000a8793
00700293
fa88cae3
01412f83
02412f03
00040613
000c8e93
000d8c93
00078d93
000a0793
00098413
00090a13
00068993
00078913
000b8693
000d0b93
00060d13
01a989b3
00170713
018da023
01ada223
05312423
04e12223
00700613
008d8d93
eae65663
04010613
000a0593
000b0513
03d12623
02d12423
03e12223
01f12a23
af8ff0ef
f6051263
04812983
04412703
02c12e83
02812683
02412f03
01412f83
000a8d93
e68ff06f
04010613
000a0593
000b0513
03d12423
02d12223
01e12a23
ab8ff0ef
f2051263
04812983
04412703
02812e83
02412683
01412f03
000a8d93
e90ff06f
01000693
04412703
0796d063
01000d13
00700413
00c0006f
ff0c8c93
059d5663
01098993
00170713
0187a023
01a7a223
05312423
04e12223
00878793
fce45ee3
04010613
000a0593
000b0513
a48ff0ef
ea051a63
ff0c8c93
04812983
04412703
000a8793
fb9d4ee3
019989b3
00170713
0187a023
0197a223
05312423
04e12223
00700793
e4e7d863
04010613
000a0593
000b0513
a00ff0ef
e6051663
04812983
e34ff06f
00040a13
e5cff06f
840e9ee3
000d0693
00000e93
00000c93
0f010413
85dff06f
2006f613
38061c63
41f75b93
00070c93
000b8613
809ff06f
00812783
010d7693
0007a703
00478793
00f12423
02069463
040d7693
00068c63
01071c93
010cdc93
00000b93
00100613
861ff06f
200d7693
32069e63
00070c93
00000b93
00100613
849ff06f
00812783
0106f613
0007a703
00478793
00f12423
02061263
0406f613
00060a63
01071c93
010cdc93
00000b93
925ff06f
2006f613
30061c63
00070c93
00000b93
911ff06f
400d7793
00000713
03312223
03412423
03212623
000c8993
000b8a13
01812903
0f010413
01d12a23
00078c93
00070b93
0240006f
00a00613
00000693
00098513
000a0593
511000ef
240a0c63
00050993
00058a13
00a00613
00000693
00098513
000a0593
2b0010ef
03050513
fea40fa3
001b8b93
fff40413
fa0c8ee3
00094683
fb769ae3
0ff00793
fafb86e3
140a1e63
00900793
1537ea63
0f010793
01212c23
01412e83
02412983
02812a03
02c12903
40878cb3
000d0693
ef8ff06f
01812783
00094603
b4078e63
0007c783
b4078a63
40046413
b4cff06f
0007a703
00412783
00c12423
41f7d693
00f72023
00d72223
aa4ff06f
00040d13
fc0ff06f
00025737
ea470793
00040693
00f12823
0206f713
06070263
00812783
00778793
ff87f793
0007ac83
0047ab83
00878793
00f12423
0016f593
00058e63
017ce5b3
00058a63
03000593
02b10e23
02c10ea3
0026e693
bff6fd13
00200613
ea8ff06f
00025737
eb870793
00040693
00f12823
0206f713
fa0712e3
00812783
0106f593
0007a703
00478793
00f12423
0a059463
0406f593
08058c63
01071c93
010cdc93
00000b93
f91ff06f
00040693
f40ff06f
00040513
808e80ef
01412683
00050c93
01a12423
00000e93
decff06f
04000593
ee5e60ef
00aa2023
00aa2823
18050263
04000793
00fa2a23
960ff06f
01c12783
02012583
00000b93
40f40433
00078613
00040513
b84f30ef
00194583
00a00613
00000693
00b03833
00098513
000a0593
01090933
335000ef
e29ff06f
2006f593
0a059663
00070c93
00000b93
ef9ff06f
00090a13
b58ff06f
00194603
02046413
00190913
9d0ff06f
00194603
20046413
00190913
9c0ff06f
00812783
0007a703
00412783
00c12423
00f72023
91cff06f
00600713
000e8c93
01d77463
00600c93
00025337
000c8b93
01a12423
ecc30413
9f8ff06f
00900793
db37e4e3
df1ff06f
04010613
000a0593
000b0513
e71fe0ef
adcff06f
00812783
00c12423
0007a703
00412783
00f71023
8c0ff06f
0ff77c93
00000b93
e51ff06f
0ff77c93
00000b93
00100613
d10ff06f
01871c93
418cdc93
41fcdb93
000b8613
c70ff06f
0ff77c93
00000b93
dfcff06f
000e8c93
01a12423
00000e93
c90ff06f
00068d13
c74ff06f
fff00793
00f12223
a70ff06f
00812783
0007ae83
00478793
000ed463
fff00e93
00194603
00f12423
00070913
8c8ff06f
00c00793
00fb2023
fff00793
00f12223
a38ff06f
fe010113
00812c23
00912a23
040017b7
00112e23
9307a783
00050413
00068493
02058263
000780e7
fff00793
02f50663
01c12083
01812403
01412483
02010113
00008067
00000613
00410593
000780e7
fff00793
fcf51ee3
0004a023
08a00793
01c12083
00f42023
01812403
01412483
02010113
00008067
fe010113
040017b7
00812c23
00912a23
00112e23
9e47a483
040017b7
9307a783
00060413
02050a63
00058613
00040693
00050593
00048513
000780e7
fff00793
02f50a63
01c12083
01812403
01412483
02010113
00008067
00060693
00410593
00000613
00048513
000780e7
fff00793
fcf51ae3
00042023
01c12083
01812403
08a00793
00f4a023
01412483
02010113
00008067
ff010113
00600513
00112623
368000ef
00100513
6e0000ef
000257b7
0d07a703
14872783
04078c63
0047a703
01f00813
06e84e63
00271813
02050663
01078333
08c32423
1887a883
00100613
00e61633
00c8e8b3
1917a423
10d32423
00200693
02d50463
00170713
00e7a223
010787b3
00b7a423
00000513
00008067
14c70793
14f72423
fa5ff06f
18c7a683
00170713
00e7a223
00c6e6b3
18d7a623
010787b3
00b7a423
00000513
00008067
fff00513
00008067
2dc52783
00078663
00000513
00008067
ff010113
08000593
00812423
00112623
00050413
b5de60ef
2ca42e23
02050463
08050793
00052023
00450513
fef51ce3
00000513
00c12083
00812403
01010113
00008067
fff00513
fedff06f
fe010113
00912a23
00112e23
00812c23
01f00793
00050493
02b7ea63
2dc52703
00058413
04070463
00241413
00870733
00072503
00c72023
01c12083
01812403
01412483
02010113
00008067
01c12083
01812403
01600793
00f52023
01412483
fff00513
02010113
00008067
08000593
00c12623
ab1e60ef
2ca4ae23
00050713
02050063
00c12603
00050793
08050693
0007a023
00478793
fed79ce3
f8dff06f
fff00513
f95ff06f
ff010113
00912223
00112623
00812423
01f00793
00050493
0ab7ea63
2dc52783
00058413
04078463
00259713
00e787b3
0007a703
02070c63
00100693
06d70c63
fff00693
04d70863
00058513
0007a023
000700e7
00000513
00c12083
00812403
00412483
01010113
00008067
00048513
484000ef
00040613
00812403
00c12083
00050593
00048513
00412483
01010113
3fc0006f
00c12083
00812403
01600793
00f52023
00412483
00100513
01010113
00008067
00c12083
00812403
00412483
00000513
01010113
00008067
01600793
00f52023
fff00513
f81ff06f
01f00793
0cb7ea63
2dc52703
ff010113
00812423
00912223
00112623
00058413
00050493
06070063
00241793
00f70733
00072783
02078c63
fff00693
08d78663
00100693
06d78663
00040513
00072023
000780e7
00000513
00c12083
00812403
00412483
01010113
00008067
00c12083
00812403
00412483
00100513
01010113
00008067
08000593
919e60ef
2ca4ae23
00050713
02050e63
00050793
08050693
0007a023
00478793
fed79ce3
f7dff06f
00c12083
00812403
00412483
00300513
01010113
00008067
00200513
f8dff06f
fff00513
f85ff06f
fff00513
00008067
ff010113
00912223
04001737
00112623
00812423
01f00793
9e472483
0aa7e863
2dc4a783
00050413
04078263
00251713
00e787b3
0007a703
02070a63
00100693
06d70a63
fff00693
04d70663
0007a023
000700e7
00000513
00c12083
00812403
00412483
01010113
00008067
00048513
2c8000ef
00040613
00812403
00c12083
00050593
00048513
00412483
01010113
2400006f
00c12083
00812403
01600793
00f4a023
00100513
00412483
01010113
00008067
00c12083
00812403
00412483
00000513
01010113
00008067
01600793
00f4a023
fff00513
f81ff06f
ff010113
01212023
04001737
00112623
00812423
00912223
01f00793
9e472903
02a7ee63
00050413
2dc92503
00058493
04050863
00241413
008507b3
0007a503
0097a023
00c12083
00812403
00412483
00012903
01010113
00008067
00c12083
00812403
01600793
00f92023
00412483
00012903
fff00513
01010113
00008067
08000593
00090513
f5ce60ef
2ca92e23
00050e63
00050793
08050713
0007a023
00478793
fee79ce3
f8dff06f
fff00513
f95ff06f
ff010113
040017b7
00812423
9e47a403
00112623
2dc42783
00078c63
00000513
00c12083
00812403
01010113
00008067
08000593
00040513
ef8e60ef
2ca42e23
00050c63
08050793
00052023
00450513
fef51ce3
fc9ff06f
fff00513
fc5ff06f
ff010113
00912223
04001737
00112623
00812423
01f00793
9e472483
0aa7ee63
2dc4a703
00050413
06070063
00241793
00f70733
00072783
02078c63
fff00693
08d78863
00100693
06d78863
00040513
00072023
000780e7
00000513
00c12083
00812403
00412483
01010113
00008067
00c12083
00812403
00412483
00100513
01010113
00008067
08000593
00048513
e40e60ef
2ca4ae23
00050713
02050e63
00050793
08050693
0007a023
00478793
fed79ce3
f79ff06f
00c12083
00812403
00412483
00300513
01010113
00008067
00200513
f89ff06f
fff00513
f81ff06f
ff010113
00058713
00812423
00912223
00050413
042594b7
00060593
00070513
00112623
b404a823
160000ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
b504a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
0d80006f
ff010113
00112623
00812423
03900893
00000073
00050413
00054c63
00c12083
00040513
00812403
01010113
00008067
40800433
f4dfa0ef
00852023
fff00413
fddff06f
05d00893
00000073
00054463
0000006f
ff010113
00812423
00050413
00112623
40800433
f19fa0ef
00852023
0000006f
f7010113
08912223
08112623
00058493
08812423
05000893
00010593
00000073
00050413
02054463
00048513
00010593
0e0000ef
08c12083
00040513
08812403
08412483
09010113
00008067
40800433
ebdfa0ef
00852023
fff00413
fcdff06f
00100513
00008067
f9010113
00810593
06112623
f8dff0ef
fff00793
00f50e63
00c12503
06c12083
00d55513
00157513
07010113
00008067
06c12083
00000513
07010113
00008067
ff010113
00112623
e5dfa0ef
00c12083
01600793
00f52023
fff00513
01010113
00008067
ff010113
00112623
00812423
03e00893
00000073
00050413
00054c63
00c12083
00040513
00812403
01010113
00008067
40800433
e0dfa0ef
00852023
fff00413
fddff06f
ff010113
0145a383
0185a283
01c5af83
0205af03
0305ae83
0405ae03
0385a303
0485a803
04c5a883
0585a603
00812623
00912423
0105a403
0085a483
01212223
0005a903
05c5a683
0685a703
06c5a783
01251023
00951123
00852223
00751423
00551523
01f51623
01e51723
01d52823
05c52623
04652423
01052c23
01152e23
02c52423
02d52623
00c12403
02e52c23
02f52e23
00812483
00412903
01010113
00008067
fd010113
01312e23
02112623
02812423
02912223
03212023
01412c23
01512a23
01612823
01712623
01812423
01912223
00050993
38069463
000257b7
00060a13
00050493
c0878793
12c5f863
00010737
00058913
10e67863
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
02000693
00e787b3
40f68733
00f68c63
00e59933
00f9d7b3
00e61a33
0127e933
00e994b3
010a5a93
000a8593
00090513
010a1b13
c8ce50ef
010b5b13
00050593
00050993
000b0513
c4ce50ef
00050413
000a8593
00090513
cb0e50ef
01051513
0104d713
00a76733
00098913
00877e63
01470733
fff98913
01476863
00877663
ffe98913
01470733
40870433
000a8593
00040513
c2ce50ef
00050593
00050993
000b0513
bf0e50ef
00050b13
000a8593
00040513
c54e50ef
01049713
01051513
01075713
00a76733
00098693
01677c63
00ea0733
fff98693
01476663
01677463
ffe98693
01091793
00d7e7b3
00000913
1200006f
010006b7
01000713
eed66ce3
01800713
ef1ff06f
00061463
00100073
00010737
12e67c63
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
02000693
00e787b3
40f68733
12f69263
40c589b3
00100913
010a5b13
000b0593
00098513
010a1b93
b68e50ef
010bdb93
00050593
00050c13
000b8513
b28e50ef
00050a93
000b0593
00098513
b8ce50ef
01051513
0104d713
00a76733
000c0993
01577e63
01470733
fffc0993
01476863
01577663
ffec0993
01470733
41570433
000b0593
00040513
b08e50ef
00050593
00050a93
000b8513
acce50ef
00050b93
000b0593
00040513
b30e50ef
01049713
01051513
01075713
00a76733
000a8693
01777c63
00ea0733
fffa8693
01476663
01777463
ffea8693
01099793
00d7e7b3
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00090593
00078513
02012903
03010113
00008067
010006b7
01000713
ecd668e3
01800713
ec9ff06f
00e61a33
00f5d933
010a5b93
00e595b3
00f9d7b3
00b7eab3
00e994b3
000b8593
00090513
010a1993
a38e50ef
0109d993
00050593
00050b13
00098513
9f8e50ef
00050413
000b8593
00090513
a5ce50ef
01051513
010ad713
00a76733
000b0913
00877e63
01470733
fffb0913
01476863
00877663
ffeb0913
01470733
40870433
000b8593
00040513
9d8e50ef
00050593
00050b13
00098513
99ce50ef
00050993
000b8593
00040513
a00e50ef
010a9793
01051513
0107d793
00a7e7b3
000b0713
0137fe63
014787b3
fffb0713
0147e863
0137f663
ffeb0713
014787b3
01091913
413789b3
00e96933
e01ff06f
1ed5ec63
000107b7
04f6f463
1006b513
00154513
00351513
000257b7
00a6d733
c0878793
00e787b3
0007c703
02000793
00a70733
40e78933
02e79663
00100793
e8b6e2e3
00c9b7b3
0017c793
e79ff06f
010007b7
01000513
fcf6e0e3
01800513
fb9ff06f
012696b3
00e65b33
00db6b33
00e5da33
010b5c13
00e9d733
012595b3
00b76ab3
000a0513
000c0593
010b1b93
012614b3
010bdb93
8dce50ef
00050593
00050c93
000b8513
8a0e50ef
00050413
000c0593
000a0513
904e50ef
01051513
010ad693
00a6e6b3
000c8a13
0086fe63
016686b3
fffc8a13
0166e863
0086f663
ffec8a13
016686b3
40868433
000c0593
00040513
880e50ef
00050593
00050c93
000b8513
844e50ef
00050b93
000c0593
00040513
8a8e50ef
010a9713
01051513
01075713
00a76733
000c8693
01777e63
01670733
fffc8693
01676863
01777663
ffec8693
01670733
010a1793
00010e37
00d7e7b3
fffe0313
41770833
0067f733
0064f333
0107de93
0104d493
00070513
00030593
fd5e40ef
00050893
00048593
00070513
fc5e40ef
00050713
00030593
000e8513
fb5e40ef
00050313
00048593
000e8513
fa5e40ef
00670733
0108d693
00d70733
00677463
01c50533
01075693
00a686b3
02d86663
bcd81ce3
00010637
fff60613
00c77733
01071713
00c8f8b3
012996b3
01170733
00000913
cce6fce3
fff78793
badff06f
00000913
00000793
cc5ff06f
fd010113
02812423
02912223
02112623
03212023
01312e23
01412c23
01512a23
01612823
01712623
01812423
01912223
01a12023
00050413
00058493
24069c63
000257b7
00060a13
c0878793
12c5fe63
00010737
12e67063
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
00e787b3
02000713
40f70933
00f70c63
012595b3
00f557b3
01261a33
00b7e4b3
01251433
010a5a93
000a8593
010a1b13
00048513
ecde40ef
010b5b13
000b0593
e95e40ef
00050993
000a8593
00048513
ef9e40ef
01051513
01045793
00a7e7b3
0137fa63
014787b3
0147e663
0137f463
014787b3
413784b3
000a8593
00048513
e81e40ef
000b0593
e4de40ef
00050993
000a8593
00048513
eb1e40ef
01041413
01051513
01045413
00a46433
01347a63
01440433
01446663
01347463
01440433
41340433
01245533
00000593
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00012d03
03010113
00008067
010006b7
01000713
eed664e3
01800713
ee1ff06f
00061463
00100073
00010737
0ee67663
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
40c584b3
00e787b3
02000713
40f70933
ecf70ae3
01261a33
00f5dbb3
010a5b13
00f557b3
012595b3
00b7e9b3
01251433
000b0593
010a1a93
000b8513
d85e40ef
010ada93
000a8593
d4de40ef
00050493
000b0593
000b8513
db1e40ef
01051513
0109d713
00a76733
00977a63
01470733
01476663
00977463
01470733
409704b3
000b0593
00048513
d39e40ef
000a8593
d05e40ef
00050a93
000b0593
00048513
d69e40ef
01099793
01051513
0107d793
00a7e7b3
0157fa63
014787b3
0147e663
0157f463
014787b3
415784b3
e19ff06f
010006b7
01000713
f0d66ee3
01800713
f15ff06f
ead5e4e3
000107b7
04f6fe63
1006b793
0017c793
00379793
00025737
00f6d833
c0870713
01070733
00074983
00f989b3
02000793
41378933
05379063
00b6e463
00c56c63
40c50633
40d586b3
00c535b3
40b684b3
00060413
00040513
00048593
e49ff06f
01000737
01000793
fae6e6e3
01800793
fa5ff06f
012696b3
01365b33
00db6b33
0135d4b3
01355a33
012595b3
010b5c93
00ba6a33
01251ab3
000c8593
00048513
010b1c13
01261bb3
010c5c13
c2de40ef
00050593
00050d13
000c0513
bf1e40ef
00050413
000c8593
00048513
c55e40ef
01051513
010a5793
00a7e7b3
000d0493
0087fe63
016787b3
fffd0493
0167e863
0087f663
ffed0493
016787b3
40878433
000c8593
00040513
bd1e40ef
00050593
00050d13
000c0513
b95e40ef
000c8593
00050c13
00040513
bf9e40ef
010a1593
01051513
0105d593
00a5e5b3
000d0793
0185fe63
016585b3
fffd0793
0165e863
0185f663
ffed0793
016585b3
00010eb7
01049493
00f4e4b3
fffe8793
00f4f8b3
00fbf7b3
41858733
0104d493
010bde13
00088513
00078593
b25e40ef
00050813
000e0593
00088513
b15e40ef
00050893
00078593
00048513
b05e40ef
00050313
000e0593
00048513
af5e40ef
01085793
006888b3
011787b3
00050613
0067f463
01d50633
0107d693
00c686b3
00010637
fff60613
00c7f7b3
01079793
00c87833
010787b3
00d76663
00d71e63
00fafc63
41778633
00c7b7b3
016787b3
40f686b3
00060793
40fa87b3
00fabab3
40d705b3
415585b3
013599b3
0127d7b3
00f9e533
0125d5b3
c71ff06f
00100837
fff80813
fe010113
00b878b3
0145d713
01d55793
00d87833
00812c23
7ff77413
00389713
0146d893
00381813
00912a23
00e7e7b3
7ff8f893
01d65713
00112e23
01212823
01312623
01f5d493
01f6d693
01076733
00351513
00361613
41140833
2cd49863
13005063
04089063
00c766b3
70068e63
fff80593
02059063
00c50633
00e78733
00a637b3
00f707b3
00060513
00100413
0700006f
7ff00693
02d81063
7ff00413
2140006f
7ff00693
20d40663
008006b7
00d76733
00080593
03800693
0ab6cc63
01f00693
06b6ce63
02000813
40b80833
010716b3
00b658b3
01061833
0116e6b3
01003833
0106e6b3
00b755b3
00a686b3
00f585b3
00a6b7b3
00f587b3
00068513
00800737
00e7f733
1a070663
00140413
7ff00713
5ce40a63
ff800737
fff70713
00e7f7b3
00155713
00157513
00a76733
01f79513
00e56533
0017d793
1780006f
fe058693
02000893
00d756b3
00000813
01158863
04000813
40b80833
01071833
00c86833
01003833
0106e6b3
00000593
f7dff06f
00c766b3
00d036b3
ff1ff06f
0e080263
408885b3
02041e63
00a7e6b3
52068c63
fff58693
00069c63
00c50533
00e78733
00c53633
00c707b3
ee1ff06f
7ff00813
03059263
00070793
00060513
eddff06f
7ff00693
fed888e3
008006b7
00d7e7b3
00058693
03800593
06d5ce63
01f00593
04d5c063
02000813
40d80833
010795b3
00d55333
01051833
0065e5b3
01003833
0105e5b3
00d7d6b3
00c58533
00e686b3
00c53633
00c687b3
00088413
ee1ff06f
fe068593
02000313
00b7d5b3
00000813
00668863
04000813
40d80833
01079833
00a86833
01003833
0105e5b3
00000693
fb9ff06f
00a7e5b3
00b035b3
ff1ff06f
00140693
7fe6f593
08059863
00a7e6b3
06041463
46068063
00c766b3
02068a63
00c50633
00e78733
00a637b3
00f707b3
00800737
00e7f733
00060513
00070a63
ff800737
fff70713
00e7f7b3
00100413
00757713
42070c63
00f57713
00400693
42d70663
00450713
00a73533
00a787b3
00070513
4180006f
ec068ee3
00c76733
da070ce3
00000493
004007b7
00000513
7ff00413
3f80006f
7ff00593
3eb68263
00c50633
00a63533
00e78733
00a70733
01f71513
00165613
00c56533
00175793
00068413
f8dff06f
0f005c63
08089e63
00c766b3
44068863
fff80593
02059063
40c50633
40e78733
00c537b3
40f707b3
00060513
00100413
0540006f
7ff00693
d2d80ce3
03800693
0ab6c663
01f00693
06b6c863
02000813
40b80833
010716b3
00b658b3
01061833
0116e6b3
01003833
0106e6b3
00b755b3
40d506b3
40b785b3
00d537b3
40f587b3
00068513
00800937
0127f733
ee070ee3
fff90913
0127f933
00050993
2140006f
7ff00693
eed402e3
008006b7
00d76733
00080593
f89ff06f
fe058693
02000893
00d756b3
00000813
01158863
04000813
40b80833
01071833
00c86833
01003833
0106e6b3
00000593
f89ff06f
00c766b3
00d036b3
ff1ff06f
0e080863
40888833
04041263
00a7e5b3
34058e63
fff80593
00059e63
40a60533
40f70733
00a63633
40c707b3
00068493
f05ff06f
7ff00313
02681463
00070793
00060513
7ff00413
0d00006f
7ff00593
feb886e3
008005b7
00b7e7b3
00080593
03800813
08b84063
01f00813
04b84263
02000313
40b30333
00b55e33
00679833
00651333
01c86833
00603333
00686533
00b7d5b3
40a60533
40b705b3
00a63633
40c587b3
00088413
00068493
ee1ff06f
fe058813
02000e13
0107d833
00000313
01c58863
04000313
40b30333
00679333
00a36333
00603333
00686533
00000593
fb5ff06f
00a7e533
00a03533
ff1ff06f
00140593
7fe5f593
08059863
00a7e833
00c765b3
06041263
00081c63
26058863
00070793
00060513
00068493
d75ff06f
d60588e3
40c50833
010538b3
40e785b3
411585b3
008008b7
0115f8b3
00088c63
40a60533
40f70733
00a63633
40c707b3
fc9ff06f
00b86533
22050a63
00058793
00080513
d2dff06f
00081c63
22058463
00070793
00060513
00068493
afdff06f
ae058ce3
d41ff06f
40c509b3
013535b3
40e78933
40b90933
008005b7
00b975b3
08058463
40a609b3
40f70933
01363633
40c90933
00068493
08090263
00090513
76c050ef
ff850713
01f00793
08e7c063
02000793
40e787b3
00e91933
00f9d7b3
0127e7b3
00e99533
0a874463
40870733
00170613
01f00693
06c6c263
02000713
40c70733
00e796b3
00c555b3
00e51733
00b6e6b3
00e03733
00e6e533
00c7d7b3
00000413
c6dff06f
0129e533
f80516e3
00000793
00000413
14c0006f
00098513
6ec050ef
02050513
f7dff06f
fd850793
00f997b3
00000513
f91ff06f
fe170713
02000593
00e7d733
00000693
00b60863
04000693
40c686b3
00d796b3
00d566b3
00d036b3
00d76533
00000793
f95ff06f
40e40433
ff800737
fff70713
00e7f7b3
bf1ff06f
00070793
00060513
00058413
be1ff06f
00070793
00060513
bd5ff06f
7ff00413
00000793
00000513
00800737
00e7f733
00070e63
00140413
7ff00713
0ce40263
ff800737
fff70713
00e7f7b3
01d79693
00355513
7ff00713
00a6e6b3
0037d793
00e41e63
00f6e6b3
00000793
00068863
000807b7
00000693
00000493
01441713
7ff00637
00c79793
01c12083
01812403
00c77733
00c7d793
01f49493
00f767b3
0097e733
01012903
01412483
00c12983
00068513
00070593
02010113
00008067
00080413
b29ff06f
00070793
00060513
00080413
da1ff06f
00000793
00000513
00000493
f45ff06f
00000793
ff5ff06f
00000513
00000493
004007b7
b31ff06f
00000793
00000513
f45ff06f
fb010113
05212023
0145d913
04912223
03312e23
03412c23
03512a23
03612823
00c59493
04112623
04812423
03712623
03812423
03912223
03a12023
01b12e23
7ff97913
00050993
00060b13
00068a93
00c4d493
01f5da13
0a090063
7ff00793
0ef90e63
01d55c93
00349493
009cecb3
008007b7
00fcecb3
00351413
c0190913
00000b93
014ad793
00ca9993
7ff7f793
00c9d993
01fada93
10078063
7ff00713
16e78063
00399993
01db5713
01376733
008009b7
013769b3
003b1813
c0178793
00000713
40f90933
002b9793
00e7e7b3
fff78793
00e00693
015a44b3
14f6ee63
000256b7
00279793
bcc68693
00d787b3
0007a783
00078067
00a4ecb3
060c8e63
04048063
00048513
474050ef
ff550793
01c00713
02f74c63
01d00c93
ff850413
40fc8cb3
008494b3
0199dcb3
009cecb3
00899433
c0d00913
40a90933
f45ff06f
43c050ef
02050513
fc5ff06f
fd850c93
01999cb3
00000413
fddff06f
00a4ecb3
020c8463
00050413
00048c93
7ff00913
00300b93
f11ff06f
00000413
00000913
00100b93
f01ff06f
00000413
7ff00913
00200b93
ef1ff06f
0169e833
06080e63
04098063
00098513
3d4050ef
ff550713
01c00793
02e7ce63
01d00793
ff850813
40e787b3
010999b3
00fb57b3
0137e9b3
010b1833
c0d00793
40a787b3
ee5ff06f
000b0513
398050ef
02050513
fc1ff06f
fd850993
013b19b3
00000813
fd9ff06f
0169e833
02080263
000b0813
7ff00793
00300713
eb1ff06f
00000993
00000793
00100713
ea1ff06f
00000993
7ff00793
00200713
e91ff06f
0199e663
453c9a63
45046863
01fc9713
00145793
01f41d93
001cdc93
00f76433
01885a93
00899b93
017aeab3
010bdb93
000b8593
010a9c13
000c8513
00881b13
010c5c13
848e40ef
00050593
00050d13
000c0513
80ce40ef
00050993
000b8593
000c8513
870e40ef
01051513
01045713
00a76733
000d0a13
01377e63
01570733
fffd0a13
01576863
01377663
ffed0a13
01570733
413709b3
000b8593
00098513
fede30ef
00050593
00050d13
000c0513
fb1e30ef
00050c93
000b8593
00098513
814e40ef
01041413
01051513
01045413
00a46433
000d0793
01947e63
01540433
fffd0793
01546863
01947663
ffed0793
01540433
010a1713
00010337
00f76733
41940433
fff30c93
019777b3
019b7cb3
01075e13
010b5d13
00078513
000c8593
f41e30ef
00050813
000d0593
00078513
f31e30ef
00050793
000c8593
000e0513
f21e30ef
00050893
000d0593
000e0513
f11e30ef
01085a13
011787b3
00fa0a33
00050693
011a7463
006506b3
010a5793
00d787b3
000106b7
fff68693
00da7a33
010a1a13
00d87833
010a0a33
00f46863
00070993
04f41463
054df263
016d8db3
016db6b3
015686b3
00d40433
fff70993
008ae663
028a9463
036de263
00f46663
00879e63
014dfc63
016d8db3
ffe70993
016db733
01570733
00e40433
414d8a33
40f40433
014db7b3
40f40433
fff00813
1a8a8263
000b8593
00040513
e91e30ef
00050593
00a12623
000c0513
e55e30ef
00a12423
000b8593
00040513
eb9e30ef
00c12683
00812783
01051513
010a5713
00a76733
00068d93
00f77e63
01570733
fff68d93
01576863
00f77663
ffe68d93
01570733
40f70433
000b8593
00040513
e2de30ef
00050593
00a12423
000c0513
df1e30ef
00050c13
000b8593
00040513
e55e30ef
00812783
010a1713
01051513
01075713
00a76733
00078693
01877e63
01570733
fff78693
01576863
01877663
ffe78693
01570733
010d9793
00d7e7b3
01079813
01085813
41870733
0107de13
00080513
000c8593
d89e30ef
00050893
000d0593
00080513
d79e30ef
00050813
000c8593
000e0513
d69e30ef
00050313
000d0593
000e0513
d59e30ef
0108d693
00680833
010686b3
00050593
0066f663
00010637
00c505b3
0106d613
00b60633
000105b7
fff58593
00b6f6b3
01069693
00b8f8b3
011686b3
00c76863
24c71a63
00078813
04068063
00ea8733
fff78813
03576463
00c76663
22c71a63
02db7063
ffe78813
001b1793
0167bb33
015b0b33
01670733
00078b13
00c71463
00db0463
00186813
3ff90793
12f05063
00787713
02070063
00f87713
00400693
00d70a63
00480713
01073833
010989b3
00070813
01000737
00e9f733
00070a63
ff0007b7
fff78793
00f9f9b3
40090793
7fe00713
0af74663
00385813
01d99713
01076733
0039d593
7ff006b7
01479793
00c59593
04c12083
04812403
00d7f7b3
00c5d593
00b7e7b3
01f49493
0097e6b3
04012903
04412483
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
00070513
00068593
05010113
00008067
fff90913
00000d93
bc1ff06f
000a0493
000c8993
00040813
000b8713
00300793
10f70063
00100793
0ef70663
00200793
f0f716e3
00000593
00000713
7ff00793
f5dff06f
000a8493
fd5ff06f
000809b7
00000813
00000493
00300713
fc1ff06f
00100593
40f585b3
03800713
0ab74463
01f00713
06b74663
41e90913
012997b3
00b85733
01281933
00e7e7b3
01203933
0127e7b3
00b9d5b3
0077f713
02070063
00f7f713
00400693
00d70a63
00478713
00f737b3
00f585b3
00070793
00800737
00e5f733
06071863
01d59713
0037d793
00f76733
0035d593
00000793
ec1ff06f
fe100713
40f707b3
02000693
00f9d7b3
00000713
00d58663
43e90713
00e99733
01076733
00e03733
00e7e7b3
00000593
f89ff06f
00000593
00000713
fbdff06f
000805b7
00000713
7ff00793
00000493
e6dff06f
00000593
00000713
00100793
e5dff06f
00080793
00078813
dedff06f
0145d713
001007b7
fff78793
0146d813
00050313
00050e93
7ff77713
7ff00513
00b7f8b3
00060f13
00d7f7b3
01f5d593
7ff87813
01f6d693
00a71c63
0068ee33
00100513
000e1463
00e80663
00008067
00a81863
00c7e633
00100513
fe0618e3
00100513
ff0714e3
fef892e3
ffee90e3
00d58a63
fc071ce3
0068e8b3
01103533
00008067
00000513
00008067
00100737
fff70713
0145d813
00b778b3
00050793
00050313
7ff87813
01f5d513
7ff00e93
0146d593
00d77733
00060e13
7ff5f593
01f6d693
01d81a63
00f8eeb3
080e8a63
ffe00513
00008067
01d59663
00c76eb3
fe0e98e3
08081063
00f8e7b3
0017b793
00059663
00c76633
04060c63
00079c63
00d51463
0305d063
04050063
fff00513
00008067
fff00513
00068a63
00068513
00008067
00b85663
fe0502e3
00008067
fd176ce3
02e89263
fc6e68e3
ffc366e3
00000513
00008067
00100513
00008067
fe0798e3
fb5ff06f
fce8e8e3
fe5ff06f
f7058ee3
f8059ee3
00000793
f89ff06f
00100737
fff70713
0145d813
00b778b3
00050793
00050313
7ff87813
01f5d513
7ff00e93
0146d593
00d77733
00060e13
7ff5f593
01f6d693
01d81a63
00f8eeb3
080e8a63
00200513
00008067
01d59663
00c76eb3
fe0e98e3
08081063
00f8e7b3
0017b793
00059663
00c76633
04060c63
00079c63
00d51463
0305d063
04050063
fff00513
00008067
fff00513
00068a63
00068513
00008067
00b85663
fe0502e3
00008067
fd176ce3
02e89263
fc6e68e3
ffc366e3
00000513
00008067
00100513
00008067
fe0798e3
fb5ff06f
fce8e8e3
fe5ff06f
f7058ee3
f8059ee3
00000793
f89ff06f
fd010113
01312e23
0145d993
02812423
02912223
01412c23
01512a23
01712623
00c59493
02112623
03212023
01612823
7ff9f993
00050413
00060b93
00068a13
00c4d493
01f5da93
3c098863
7ff00793
42f98663
00349493
01d55793
0097e7b3
008004b7
0097e4b3
00351913
c0198993
00000b13
014a5713
00ca1413
7ff77713
00c45413
01fa5a13
42070663
7ff00793
48f70663
00341413
01dbd793
0087e7b3
00800437
0087e433
c0170713
003b9793
00000613
00e989b3
002b1713
00c76733
00a00693
014ac833
00198893
4ce6c863
00200693
48e6c063
fff70713
00100693
48e6fc63
00010a37
fffa0393
0107d293
00797e33
0077f7b3
01095f93
000e0513
00078593
f60e30ef
00050e93
00028593
000e0513
f50e30ef
00050713
00078593
000f8513
f40e30ef
00050913
00028593
000f8513
f30e30ef
010ed313
01270733
00e30333
00050f13
01237463
01450f33
01035913
00737333
007efeb3
01031313
007473b3
01d30333
01045a13
000e0513
00038593
ef0e30ef
00050e93
000a0593
000e0513
ee0e30ef
00050e13
00038593
000f8513
ed0e30ef
00050413
000a0593
000f8513
ec0e30ef
010ed713
008e0e33
01c70733
00050693
00877663
00010637
00c506b3
00010b37
fffb0e13
01075f93
01c77733
01071713
01cefeb3
01d70eb3
01c4fe33
00df8fb3
01d90933
0104da93
000e0513
00078593
e6ce30ef
00050413
00028593
000e0513
e5ce30ef
00050493
00078593
000a8513
e4ce30ef
00050b93
00028593
000a8513
e3ce30ef
01045793
017484b3
009787b3
00050713
0177f463
01650733
000104b7
fff48693
0107d293
00e282b3
00d7f733
00d47433
01071713
00870733
000e0513
00038593
df8e30ef
00050413
000a0593
000e0513
de8e30ef
00050e13
00038593
000a8513
dd8e30ef
00050393
000a0593
000a8513
dc8e30ef
01045793
007e0e33
01c78e33
00050593
007e7463
009505b3
000106b7
fff68693
00de77b3
00d47433
01079793
012f0f33
008787b3
01df3eb3
01f787b3
01d78533
00ef0f33
00ef3733
005506b3
00e68633
01f7b433
01d53533
010e5793
00e63733
00a46433
0056b6b3
00f40433
00e6e6b3
00d40433
00b40433
01765793
00941413
00f46433
009f1793
0067e7b3
00f037b3
017f5f13
00961713
01e7e7b3
00e7e7b3
01000737
00e47733
28070663
0017d713
0017f793
00f76733
01f41793
00f767b3
00145413
3ff88693
26d05a63
0077f713
02070063
00f7f713
00400613
00c70a63
00478713
00f737b3
00f40433
00070793
01000737
00e47733
00070a63
ff000737
fff70713
00e47433
40088693
7fe00713
2ed74e63
01d41713
0037d793
00f76733
00345413
7ff007b7
01469693
00c41413
00f6f6b3
00c45413
02c12083
0086e6b3
02812403
01f81813
0106e7b3
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00070513
00078593
03010113
00008067
00a4e933
06090c63
04048063
00048513
720040ef
ff550713
01c00793
02e7cc63
01d00793
ff850913
40e787b3
012494b3
00f457b3
0097e4b3
01241933
c0d00993
40a989b3
c15ff06f
6e8040ef
02050513
fc5ff06f
fd850493
009414b3
00000913
fddff06f
00a4e933
02090263
00050913
7ff00993
00300b13
be5ff06f
00000493
00000993
00100b13
bd5ff06f
00000493
7ff00993
00200b13
bc5ff06f
017467b3
06078e63
04040063
00040513
684040ef
ff550693
01c00793
02d7ce63
01d00713
ff850793
40d70733
00f41433
00ebd733
00876433
00fb97b3
c0d00713
40a70733
bb9ff06f
000b8513
648040ef
02050513
fc1ff06f
fd850413
008b9433
00000793
fd9ff06f
017467b3
02078263
000b8793
7ff00713
00300613
b85ff06f
00000413
00000713
00100613
b75ff06f
00000413
7ff00713
00200613
b65ff06f
00100693
00e696b3
5306f713
04071863
2406f593
12059463
0886f693
b6068ae3
000a0813
00200713
12e60863
00300713
10e60e63
00100713
dce61ce3
00000413
00000713
0bc0006f
00f00693
02d70063
00b00693
fcd706e3
000a8813
00048413
00090793
000b0613
fbdff06f
00080437
00000793
00000813
00300613
fb1ff06f
00098893
d8dff06f
00100613
40d60633
03800713
fac744e3
01f00713
06c74663
41e88893
01141733
00c7d6b3
011798b3
00d76733
011038b3
011767b3
00c45433
0077f713
02070063
00f7f713
00400693
00d70a63
00478713
00f737b3
00f40433
00070793
00800737
00e47733
06071e63
01d41713
0037d793
00f76733
00345413
00000693
d6dff06f
fe100713
40d70733
02000593
00e45733
00000693
00b60663
43e88893
011416b3
00f6e6b3
00d036b3
00d767b3
00000413
f89ff06f
00080437
7ff00693
00000813
d29ff06f
00080437
00000713
fedff06f
00000413
00000713
7ff00693
d0dff06f
00000413
00000713
00100693
cfdff06f
00100837
fff80813
fe010113
00b878b3
0145d713
01d55793
00d87833
00812c23
7ff77413
00389713
0146d893
00912a23
00e7e7b3
01f5d493
01d65713
00381813
00112e23
01212823
01312623
7ff8f893
7ff00593
00351513
01f6d693
01076733
00361613
00b89663
00c765b3
00059463
0016c693
41140833
2c969863
13005063
04089063
00c766b3
70068e63
fff80593
02059063
00c50633
00e78733
00a637b3
00f707b3
00060513
00100413
0700006f
7ff00693
02d81063
7ff00413
2140006f
7ff00693
20d40663
008006b7
00d76733
00080593
03800693
0ab6cc63
01f00693
06b6ce63
02000813
40b80833
010716b3
00b658b3
01061833
0116e6b3
01003833
0106e6b3
00b755b3
00a686b3
00f585b3
00a6b7b3
00f587b3
00068513
00800737
00e7f733
1a070663
00140413
7ff00713
5ce40a63
ff800737
fff70713
00e7f7b3
00155713
00157513
00a76733
01f79513
00e56533
0017d793
1780006f
fe058693
02000893
00d756b3
00000813
01158863
04000813
40b80833
01071833
00c86833
01003833
0106e6b3
00000593
f7dff06f
00c766b3
00d036b3
ff1ff06f
0e080263
408885b3
02041e63
00a7e6b3
52068c63
fff58693
00069c63
00c50533
00e78733
00c53633
00c707b3
ee1ff06f
7ff00813
03059263
00070793
00060513
eddff06f
7ff00693
fed888e3
008006b7
00d7e7b3
00058693
03800593
06d5ce63
01f00593
04d5c063
02000813
40d80833
010795b3
00d55333
01051833
0065e5b3
01003833
0105e5b3
00d7d6b3
00c58533
00e686b3
00c53633
00c687b3
00088413
ee1ff06f
fe068593
02000313
00b7d5b3
00000813
00668863
04000813
40d80833
01079833
00a86833
01003833
0105e5b3
00000693
fb9ff06f
00a7e5b3
00b035b3
ff1ff06f
00140693
7fe6f593
08059863
00a7e6b3
06041463
46068063
00c766b3
02068a63
00c50633
00e78733
00a637b3
00f707b3
00800737
00e7f733
00060513
00070a63
ff800737
fff70713
00e7f7b3
00100413
00757713
42070c63
00f57713
00400693
42d70663
00450713
00a73533
00a787b3
00070513
4180006f
ec068ee3
00c76733
da070ce3
00000493
004007b7
00000513
7ff00413
3f80006f
7ff00593
3eb68263
00c50633
00a63533
00e78733
00a70733
01f71513
00165613
00c56533
00175793
00068413
f8dff06f
0f005c63
08089e63
00c766b3
44068863
fff80593
02059063
40c50633
40e78733
00c537b3
40f707b3
00060513
00100413
0540006f
7ff00693
d2d80ce3
03800693
0ab6c663
01f00693
06b6c863
02000813
40b80833
010716b3
00b658b3
01061833
0116e6b3
01003833
0106e6b3
00b755b3
40d506b3
40b785b3
00d537b3
40f587b3
00068513
00800937
0127f733
ee070ee3
fff90913
0127f933
00050993
2140006f
7ff00693
eed402e3
008006b7
00d76733
00080593
f89ff06f
fe058693
02000893
00d756b3
00000813
01158863
04000813
40b80833
01071833
00c86833
01003833
0106e6b3
00000593
f89ff06f
00c766b3
00d036b3
ff1ff06f
0e080863
40888833
04041263
00a7e5b3
34058e63
fff80593
00059e63
40a60533
40f70733
00a63633
40c707b3
00068493
f05ff06f
7ff00313
02681463
00070793
00060513
7ff00413
0d00006f
7ff00593
feb886e3
008005b7
00b7e7b3
00080593
03800813
08b84063
01f00813
04b84263
02000313
40b30333
00b55e33
00679833
00651333
01c86833
00603333
00686533
00b7d5b3
40a60533
40b705b3
00a63633
40c587b3
00088413
00068493
ee1ff06f
fe058813
02000e13
0107d833
00000313
01c58863
04000313
40b30333
00679333
00a36333
00603333
00686533
00000593
fb5ff06f
00a7e533
00a03533
ff1ff06f
00140593
7fe5f593
08059863
00c765b3
00a7e833
06041263
00081c63
26058863
00070793
00060513
00068493
d75ff06f
d60588e3
40c50833
010538b3
40e785b3
411585b3
008008b7
0115f8b3
00088c63
40a60533
40f70733
00a63633
40c707b3
fc9ff06f
00b86533
22050a63
00058793
00080513
d2dff06f
00081c63
22058463
00070793
00060513
00068493
afdff06f
ae058ce3
d41ff06f
40c509b3
013535b3
40e78933
40b90933
008005b7
00b975b3
08058463
40a609b3
40f70933
01363633
40c90933
00068493
08090263
00090513
67d030ef
ff850713
01f00793
08e7c063
02000793
40e787b3
00e91933
00f9d7b3
0127e7b3
00e99533
0a874463
40870733
00170613
01f00693
06c6c263
02000713
40c70733
00e796b3
00c555b3
00e51733
00b6e6b3
00e03733
00e6e533
00c7d7b3
00000413
c6dff06f
0129e533
f80516e3
00000793
00000413
14c0006f
00098513
5fd030ef
02050513
f7dff06f
fd850793
00f997b3
00000513
f91ff06f
fe170713
02000593
00e7d733
00000693
00b60863
04000693
40c686b3
00d796b3
00d566b3
00d036b3
00d76533
00000793
f95ff06f
40e40433
ff800737
fff70713
00e7f7b3
bf1ff06f
00070793
00060513
00058413
be1ff06f
00070793
00060513
bd5ff06f
7ff00413
00000793
00000513
00800737
00e7f733
00070e63
00140413
7ff00713
0ce40263
ff800737
fff70713
00e7f7b3
01d79693
00355513
7ff00713
00a6e6b3
0037d793
00e41e63
00f6e6b3
00000793
00068863
000807b7
00000693
00000493
01441713
7ff00637
00c79793
01c12083
01812403
00c77733
00c7d793
01f49493
00f767b3
0097e733
01012903
01412483
00c12983
00068513
00070593
02010113
00008067
00080413
b29ff06f
00070793
00060513
00080413
da1ff06f
00000793
00000513
00000493
f45ff06f
00000793
ff5ff06f
00000513
00000493
004007b7
b31ff06f
00000793
00000513
f45ff06f
001007b7
fff78793
00b7f733
0145d593
00d7f7b3
7ff5f593
0146d693
7ff00813
7ff6f693
01059863
00a76733
00100513
00071c63
7ff00713
00000513
00e69663
00c7e7b3
00f03533
00008067
0145d713
001006b7
fff68793
7ff77713
3fe00613
00b7f7b3
01f5d593
04e65e63
41d00613
00e65a63
80000537
fff54513
00a58533
00008067
00d7e7b3
43300693
40e686b3
01f00613
02d64063
bed70713
00e797b3
00d55533
00a7e533
02058063
40a00533
00008067
41300693
40e68733
00e7d533
fe9ff06f
00000513
00008067
0145d713
00100637
00050693
fff60793
7ff77713
3fe00513
00b7f7b3
01f5d593
04e55a63
00000513
00059863
41e00593
fff00513
00e5d463
00008067
00c7e7b3
43300613
40e60633
01f00593
00c5cc63
bed70713
00e797b3
00c6d533
00a7e533
00008067
41300693
40e68733
00e7d533
00008067
00000513
00008067
ff010113
00112623
00812423
00912223
08050663
41f55793
00a7c433
40f40433
01f55493
00040513
31d030ef
41e00713
00a00793
40a70733
04a7c863
00b00793
40a787b3
01550513
00f457b3
00a41433
00048513
00c79793
00c7d793
01471713
01f51513
00f76733
00c12083
00a767b3
00040513
00812403
00412483
00078593
01010113
00008067
ff550513
00a417b3
00048513
00000413
fbdff06f
00000713
00000793
ff1ff06f
ff010113
00812423
00112623
00050413
06050263
289030ef
41e00713
00a00793
40a70733
04a7c063
00b00793
40a787b3
01550513
00f457b3
00a41433
00c12083
00040513
00c79793
00812403
01471713
00c7d793
00f766b3
00068593
01010113
00008067
ff550513
00a417b3
00000413
fcdff06f
00000793
00000713
fc1ff06f
00100737
0145d613
fff70793
7ff67613
3fe00693
00b7f7b3
0ac6da63
ff010113
00812423
00112623
43d00693
01f5d413
02c6da63
00100513
40850533
41f55713
800005b7
00a037b3
40e585b3
40a00533
40f585b3
00c12083
00812403
01010113
00008067
00e7e5b3
43200793
02c7d263
bcd60613
171030ef
fc040ee3
00a037b3
40b005b3
40f585b3
40a00533
fc9ff06f
43300793
40c787b3
01f00713
00f74e63
bed60613
00c59633
00f55533
00a66533
00f5d5b3
fc5ff06f
41300513
40c50533
00a5d533
00000593
fb1ff06f
00000513
00000593
00008067
fe010113
00112e23
00812c23
00912a23
01212823
01312623
01412423
01512223
01612023
00b567b3
1a078463
00050413
00058993
01f5d913
0005da63
00a037b3
40b009b3
40f989b3
40a00433
00098493
08098a63
00098513
0ed030ef
00050a93
43e00793
41578a33
43300793
0947cc63
00b00793
02fa8463
02a00793
0757cc63
02b00493
ff5a8793
415484b3
009454b3
00f999b3
0134e4b3
00f41433
00c49593
01c12083
014a1793
00c5d593
00040513
01812403
00b7e7b3
01f91913
0127e733
01412483
01012903
00c12983
00812a03
00412a83
00012b03
00070593
02010113
00008067
00040513
05d030ef
02050a93
f71ff06f
fd5a8593
00b414b3
00000413
f9dff06f
43600793
0547d063
00800613
41560633
00040513
00098593
7b8030ef
00050b13
00058493
00040513
00098593
038a8613
7d8030ef
00b56433
00803433
01646433
00048993
00800793
0357d063
02800713
ff8a8793
41570733
00e45733
00f999b3
013769b3
00f41433
ff8005b7
fff58593
00747793
00b9f5b3
02078063
00f47793
00400713
00e78a63
00440793
0087b433
008585b3
00078413
008007b7
00f5f7b3
00078c63
ff8007b7
fff78793
00f5f5b3
43f00793
41578a33
00345413
01d59793
0087e433
0035d493
ed1ff06f
00000493
00000413
00000a13
00000913
ebdff06f
00c52783
0005af03
0045af83
0085a283
00c5a583
00008737
0107d693
fff70713
01079813
01059e93
01f7d613
00e6f6b3
0105d793
00052883
00452303
00852e03
ff010113
01085813
010ede93
00e7f7b3
01f5d593
02e69063
0068e733
01c76733
01076733
00100513
04071a63
04d79863
0080006f
00e79c63
01ff6733
00576733
01d76733
00100513
02071a63
00100513
02d79663
03e89463
03f31263
025e1063
01d81e63
02b60063
00079a63
0068e533
01c56533
01056533
00a03533
01010113
00008067
00000513
ff5ff06f
00052f83
00452803
00852e03
00c52503
00c5a683
000087b7
01055613
fff78793
01069313
0106d713
0005a283
0045a883
0085ae83
00f67633
01051593
ff010113
0105d593
01f55513
01035313
00f77733
01f6d693
00f61e63
01f867b3
01c7e7b3
00b7e7b3
0c078863
ffe00513
0640006f
00f71a63
0112e7b3
01d7e7b3
0067e7b3
fe0794e3
0a061a63
01f867b3
01c7e7b3
00b7e7b3
0017b793
00071a63
0112ef33
01df6f33
006f6f33
060f0a63
00079c63
00a69463
02c75263
04050e63
fff00513
0100006f
fff00513
00068463
00068513
01010113
00008067
00e65663
fe051ae3
fddff06f
fcb36ae3
02659e63
fdcee6e3
03de1e63
fd08e2e3
01181463
fbf2eee3
fd186ee3
01181463
fc5feae3
00000513
fc1ff06f
00100513
fb9ff06f
fe0798e3
f99ff06f
fa65ece3
fe5ff06f
fbde68e3
fddff06f
f4c700e3
f6071ce3
00000793
f5dff06f
00052f83
00452803
00852e03
00c52503
00c5a683
000087b7
01055613
fff78793
01069313
0106d713
0005a283
0045a883
0085ae83
00f67633
01051593
ff010113
0105d593
01f55513
01035313
00f77733
01f6d693
00f61e63
01f867b3
01c7e7b3
00b7e7b3
0c078863
00200513
0640006f
00f71a63
0112e7b3
01d7e7b3
0067e7b3
fe0794e3
0a061a63
01f867b3
01c7e7b3
00b7e7b3
0017b793
00071a63
0112ef33
01df6f33
006f6f33
060f0a63
00079c63
00a69463
02c75263
04050e63
fff00513
0100006f
fff00513
00068463
00068513
01010113
00008067
00e65663
fe051ae3
fddff06f
fcb36ae3
02659e63
fdcee6e3
03de1e63
fd08e2e3
01181463
fbf2eee3
fd186ee3
01181463
fc5feae3
00000513
fc1ff06f
00100513
fb9ff06f
fe0798e3
f99ff06f
fa65ece3
fe5ff06f
fbde68e3
fddff06f
f4c700e3
f6071ce3
00000793
f5dff06f
f6010113
09312623
00c5a983
0005a783
0085a683
08912a23
00050493
0045a503
01099713
09412423
09512223
00c62a03
00062a83
09612023
07712e23
00862b03
00462b83
00008637
09212823
01075713
0109d913
fff60613
05312623
08112e23
08812c23
07812c23
07912a23
07a12823
07b12623
04f12023
04a12223
04d12423
00f12823
00a12a23
00d12c23
00e12e23
00c97933
01f9d993
580906e3
6ac902e3
000107b7
00f76733
00e12e23
01010613
01c10793
0007a703
ffc7a683
ffc78793
00371713
01d6d693
00d76733
00e7a223
fef612e3
01012783
00379793
00f12823
ffffc7b7
00178793
00f90933
00000c13
010a1513
00008737
010a5793
01055513
fff70713
05412623
05512023
05712223
05612423
03512023
03712223
03612423
02a12623
00e7f7b3
01fa5a13
62078ee3
00e79463
7510006f
00010737
00e56533
02a12623
02010593
02c10713
00072683
ffc72603
ffc70713
00369693
01d65613
00c6e6b3
00d72223
fee592e3
02012703
00371713
02e12023
ffffc737
00170713
00e787b3
00000693
012787b3
00f12423
00178c93
002c1793
00d7e7b3
00a00713
0149c433
00f75463
74d0006f
00200713
00f75463
6fd0006f
fff78793
00100713
00f76463
7950006f
01012283
02012f83
00010337
fff30793
00f2f833
00fff7b3
0102de93
010fd713
00080513
00078593
f39e10ef
00050e13
00070593
00080513
f29e10ef
00050813
00078593
000e8513
f19e10ef
00050893
00070593
000e8513
f09e10ef
010e5713
01180833
01070733
00050793
01177463
006507b3
01075693
00f687b3
00010337
02412e83
04f12223
fff30793
00f77733
01071713
00fe7533
00a70533
00fef833
00f2f733
04a12023
0102d893
010edf13
00070513
00080593
ea9e10ef
00050e13
000f0593
00070513
e99e10ef
00050713
00080593
00088513
e89e10ef
00050813
000f0593
00088513
e79e10ef
010e5893
01070733
00e888b3
00050a13
0108f463
00650a33
01412f03
0108d713
00f8f8b3
00fe7533
00e12623
01089893
00ff7733
00fff7b3
00a888b3
010f5393
010fd313
00070513
00078593
e29e10ef
00050813
00030593
00070513
e19e10ef
00050713
00078593
00038513
e09e10ef
00050e13
00030593
00038513
df9e10ef
01085313
01c70733
00e30333
00050793
01c37663
00010737
00e507b3
00010e37
fffe0593
01035b93
00b37333
00b87833
00bf7933
00bef3b3
01031313
00fb8bb3
01030333
010ed793
010f5813
00090513
00038593
da1e10ef
00050713
00078593
00090513
d91e10ef
00050913
00038593
00080513
d81e10ef
00050393
00078593
00080513
d71e10ef
01075813
007906b3
00d80833
00050793
00787463
01c507b3
00010e37
fffe0593
02812383
01085b13
00b87833
00b77733
01081813
00b2f933
00e80833
00b3f733
00fb0b33
0102dc13
0103da93
00090513
00070593
d19e10ef
00050793
000a8593
00090513
d09e10ef
00050993
00070593
000c0513
cf9e10ef
00050913
000a8593
000c0513
ce9e10ef
0107d713
012986b3
00d70733
01277463
01c50533
00010d37
fffd0913
01812e03
01075a93
01277733
0127f7b3
01071713
00f70733
012e77b3
012ff933
00aa8ab3
010e5d93
010fdc13
00078513
00090593
c95e10ef
00050993
000c0593
00078513
c85e10ef
00050793
00090593
000d8513
c75e10ef
00050913
000c0593
000d8513
c65e10ef
012787b3
0109d693
00d787b3
0127f463
01a50533
00010937
fff90593
04412603
0107d693
00b7f7b3
01079793
00b9f9b3
013789b3
00c12783
00c88633
011638b3
011787b3
00660633
01478a33
017a07b3
04c12223
00663633
00c78333
00a68533
0177b7b3
010306b3
00c33333
011a3a33
0067e7b3
014787b3
0106b833
016787b3
01078a33
00e686b3
00e6b733
015a08b3
00e88333
013686b3
00a30633
04d12423
0136b6b3
00d609b3
010a3a33
0167b7b3
0158b8b3
00e33333
02c12803
05312623
0147e7b3
00d9b9b3
0068e8b3
00a63633
01366633
011787b3
00c787b3
04f12823
0102da13
00b877b3
00b2f2b3
01085993
00028513
00078593
b69e10ef
00050713
00098593
00028513
b59e10ef
00050893
00078593
000a0513
b49e10ef
00050313
00098593
000a0513
b39e10ef
01075613
006888b3
01160633
00050793
00667463
012507b3
01065a13
000102b7
01c12883
00fa0a33
fff28793
00f67633
00f77733
01061613
00e60333
00f8f933
010fd713
00ffffb3
0108d993
00090513
000f8593
ae1e10ef
00050793
00070593
00090513
ad1e10ef
00050913
000f8593
00098513
ac1e10ef
00050f93
00070593
00098513
ab1e10ef
0107d693
01f90933
012686b3
00050713
01f6f463
00550733
00010fb7
ffff8613
0106d993
00c6f6b3
01069693
00c7f7b3
00cf7933
00c3f2b3
00e989b3
00f68b33
010f5713
0103da93
00090513
00028593
a5de10ef
00050793
000a8593
00090513
a4de10ef
00050913
00028593
00070513
a3de10ef
00050293
000a8593
00070513
a2de10ef
0107d713
005906b3
00d70733
00577463
01f50533
000102b7
fff28693
01075913
00d77733
00d7f7b3
00de7ab3
00deffb3
01071713
00a90933
00f70733
010e5d13
010edc13
000a8513
000f8593
9dde10ef
00050793
000c0593
000a8513
9cde10ef
00050b93
000f8593
000d0513
9bde10ef
00050a93
000c0593
000d0513
9ade10ef
0107df93
015b86b3
00df8fb3
015ff463
00550533
00010ab7
fffa8293
010fdb93
005fffb3
0057f7b3
010f9f93
00ff8fb3
04c12783
00ab8bb3
00f307b3
0067b633
05012303
016787b3
0167b6b3
006a0333
00c30d33
013d0b33
00db0c33
00e787b3
00e7b733
012c05b3
00e58533
01f787b3
04f12623
01433333
01f7b7b3
00cd3d33
01750fb3
013b3b33
00dc3c33
00ff8db3
00e53533
01a36333
018b6b33
0125b5b3
00a5e5b3
05b12823
01630333
00fdbdb3
017fbfb3
00b30333
01bfefb3
01f307b3
005e7333
0053f2b3
04f12a23
010e5913
0103d713
00030513
00028593
8cde10ef
00050793
00070593
00030513
8bde10ef
00050313
00028593
00090513
8ade10ef
00050f93
00070593
00090513
89de10ef
0107d613
01f30333
00660633
00050713
01f67463
01550733
01065993
00010fb7
00e989b3
ffff8713
00e67633
01061613
00e7f7b3
010f5a13
00ef7f33
00e87733
00f607b3
01085913
000f0513
00070593
849e10ef
00050313
00090593
000f0513
839e10ef
00050f13
00070593
000a0513
829e10ef
00050293
00090593
000a0513
819e10ef
01035693
005f0f33
01e686b3
00050713
0056f463
01f50733
000102b7
fff28613
0106d913
00c6f6b3
00c37333
01069693
00668a33
010edf13
00c8f333
00cefeb3
00e90933
00030513
0108d713
000e8593
fc4e10ef
00050f93
000f0593
00030513
fb4e10ef
00050a93
000e8593
00070513
fa4e10ef
00050313
000f0593
00070513
f94e10ef
00050713
010fdf13
006a8533
00af0f33
006f7463
00570733
010f5293
00010337
00e282b3
fff30713
00ef7f33
00efffb3
010f1f13
01ff0f33
010e5a93
00e87fb3
00ee7e33
01085b13
000e0513
000f8593
f40e10ef
00050e93
000b0593
000e0513
f30e10ef
00050713
000f8593
000a8513
f20e10ef
00050f93
000b0593
000a8513
f10e10ef
01f70733
010ed693
00d70733
01f77463
00650533
00010337
fff30593
01075f93
00b77733
00befeb3
00b8fb33
0103db93
01071713
00b3f3b3
00af8fb3
01d70733
0108de13
000b0513
00038593
ec0e10ef
00050a93
000b8593
000b0513
eb0e10ef
00050b13
00038593
000e0513
ea0e10ef
00050393
000b8593
000e0513
e90e10ef
010ade93
007b06b3
00de8eb3
007ef463
00650533
05012583
00010e37
fffe0313
00b785b3
00f5b633
05412783
014585b3
0145b6b3
00f987b3
00c78bb3
012b8a33
00da0b33
01e585b3
010ed393
006efeb3
00a383b3
006afab3
005b0533
04b12823
010e9e93
01e5b5b3
015e8eb3
00cbbbb3
00b50ab3
00db3b33
0137b7b3
012a3a33
00ea8f33
0177e7b3
00babab3
016a6a33
00553533
01556533
014787b3
00a787b3
00ef3733
01f787b3
00e785b3
01df0f33
007586b3
05e12a23
01df3f33
01e68633
00e5b5b3
04c12c23
01f7b7b3
01e63633
0076b6b3
00b7e7b3
00c6e6b3
00d787b3
04f12e23
0108df13
01085793
0068f8b3
00687833
00088513
00080593
d90e10ef
00050e93
00078593
00088513
d80e10ef
00050713
00080593
000f0513
d70e10ef
00050813
00078593
000f0513
d60e10ef
010ed793
01070733
00e787b3
00050693
0107f463
01c506b3
05812603
0067f733
05c12583
01071713
006efeb3
01d70733
00c70633
0107d793
00b787b3
00e63733
00e787b3
00d78533
04412703
04012783
04a12e23
04c12c23
00f76733
04812783
05010593
00f76733
04c12783
00d79793
00e7e7b3
04010713
00c72683
01072603
00470713
0136d693
00d61613
00c6e6b3
fed72e23
fee592e3
04812683
04012703
00f037b3
02d12c23
04412683
00e7e7b3
04c12703
02d12a23
001006b7
02e12e23
02f12823
00d77733
4e070463
01f79793
03010713
03c10593
00072683
00472603
00470713
0016d693
01f61613
00c6e6b3
fed72e23
fee592e3
03c12703
00f037b3
00175713
02e12e23
03012703
00f767b3
02f12823
000047b7
fff78793
00fc87b3
4af05863
03012703
00777693
04068463
00f77693
00400613
02c68e63
03412683
00470713
02e12823
00473713
00d706b3
02d12a23
00e6b6b3
03812703
00e68733
02e12c23
00d73733
03c12683
00d70733
02e12e23
03c12703
001006b7
00d776b3
00068e63
fff007b7
fff78793
00f77733
000047b7
02e12e23
00fc87b3
03010713
03c10593
00072683
00472603
00470713
0036d693
01d61613
00c6e6b3
fed72e23
feb712e3
000086b7
ffe68613
03c12703
3ef64463
00375713
02e12e23
01179793
0117d793
00f41413
00f46433
03012783
03c12703
04811723
00f4a023
03412783
04e11623
09c12083
00f4a223
03812783
09812403
09012903
00f4a423
04c12783
08c12983
08812a03
00f4a623
08412a83
08012b03
07c12b83
07812c03
07412c83
07012d03
06c12d83
00048513
09412483
0a010113
00008067
00a7e633
00d66633
00e66633
12060663
08070463
00070513
5d0020ef
00050413
ff440593
4055d793
01f5f593
40f00733
08058e63
00271713
00c70693
02000513
01010893
40b50533
00d886b3
40e00733
0ad89463
fff78613
00279793
01010713
05078793
00e787b3
01012703
00b71733
fae7a823
00160613
ffffc937
00261613
00000593
01010513
01190913
889e20ef
40890933
a34ff06f
00068a63
00068513
548020ef
02050413
f79ff06f
00050863
538020ef
04050413
f69ff06f
00078513
528020ef
06050413
f59ff06f
01c10693
00271713
00300613
00e685b3
0005a583
fff60613
ffc68693
00b6a223
fef656e3
fff78613
f81ff06f
0006a603
ffc6a803
00e68333
00b61633
00a85833
01066633
00c32023
ffc68693
f39ff06f
00a7e7b3
00d7e7b3
00e7e7b3
00300c13
9a079063
00200c13
998ff06f
00000913
00100c13
98cff06f
017ae7b3
0167e7b3
00a7e7b3
12078863
08050263
490020ef
00050413
ff440593
4055d793
01f5f593
40f00733
0a058063
00271713
00c70693
02000513
02010893
40b50533
00d886b3
40e00733
0ad89663
fff78613
00279793
01010713
05078793
00e787b3
02012703
00b71733
fce7a023
00160613
00261613
00000593
02010513
f50e20ef
ffffc7b7
01178793
408787b3
98cff06f
000b0a63
000b0513
408020ef
02050413
f79ff06f
000b8a63
000b8513
3f4020ef
04050413
f65ff06f
000a8513
3e4020ef
06050413
f55ff06f
02c10693
00271713
00300613
00e685b3
0005a583
fff60613
ffc68693
00b6a223
fef656e3
fff78613
f7dff06f
0006a603
ffc6a803
00e68333
00b61633
00a85833
01066633
00c32023
ffc68693
f35ff06f
017aeab3
016aeab3
00aaeab3
00300693
000a8463
8f0ff06f
00200693
8e8ff06f
00000793
00100693
8dcff06f
00100713
00f717b3
5307f713
04071663
0887f713
08071863
2407f793
00079463
8f8ff06f
000087b7
02f12e23
02012c23
02012a23
02012823
fff78793
00000413
cb9ff06f
00f00713
fce78ee3
00b00713
04e78a63
00098413
01012783
02f12823
01412783
02f12a23
01812783
02f12c23
01c12783
02f12e23
00200793
26fc0e63
00300793
fafc00e3
00100793
bafc12e3
02012e23
02012c23
02012a23
02012823
2180006f
000a0413
02012783
00068c13
02f12823
02412783
02f12a23
02812783
02f12c23
02c12783
fadff06f
00812c83
b61ff06f
02012e23
02012c23
02012a23
02012823
fff68793
c11ff06f
00100713
40f707b3
07400713
1cf74463
03010993
4057d513
00098693
00000913
00000713
04a71263
01f7f793
00251693
04079663
00300613
00098793
00000713
40a60633
00d785b3
0005a583
00170713
00478793
feb7ae23
fee656e3
00400793
40a78533
0780006f
0006a603
00170713
00468693
00c96933
fadff06f
05068713
01010613
00c70733
fd072703
02000593
40f585b3
00b71733
00e96933
00300713
00d986b3
00098893
00000813
40a70733
00468693
0ce84263
00400693
00271713
40a68533
05070713
01010693
00d70733
03c12683
00f6d7b3
fcf72823
00400a13
40aa0633
00251513
00261613
00000593
00a98533
ca8e20ef
03012703
012037b3
00e7e7b3
02f12823
0077f713
04070263
00f7f713
03470e63
03412703
00478793
02f12823
0047b793
00e78733
02e12a23
00f73733
03812783
00f707b3
02f12c23
00e7b7b3
03c12703
00e787b3
02f12e23
03c12703
000807b7
00e7f7b3
04078063
02012e23
02012c23
02012a23
02012823
00100793
a99ff06f
ffc6a603
0006a303
00180813
00f65633
00b31333
00666633
00c8a023
00488893
f19ff06f
00c98693
0009a783
0049a703
00498993
0037d793
01d71713
00e7e7b3
fef9ae23
fed992e3
03c12783
0037d793
02f12e23
00000793
a3dff06f
03412783
03012703
00f76733
03812783
00f76733
03c12783
00f76733
00000793
a0070ce3
02012e23
02012c23
02012a23
02012823
a05ff06f
000087b7
02012e23
02012c23
02012a23
02012823
fff78793
9e9ff06f
f9010113
0085a783
05312e23
00c5a983
0005a683
0045a703
05412c23
05712623
00050a13
02f12c23
00f12c23
00062883
01099793
00462503
00862583
00c62b83
06812423
0107d793
00199413
02d12823
03312e23
00d12823
06112623
06912223
07212023
05512a23
05612823
05812423
05912223
02e12a23
00e12a23
00f12e23
01145413
01f9d993
01010813
01c10693
0006a783
ffc6a703
ffc68693
00379793
01d75713
00e7e7b3
00f6a223
fed812e3
01012903
010b9793
001b9b13
00391913
0107d793
02a12a23
03712e23
02a12223
01212823
03112823
02b12c23
03112023
02b12423
02f12623
011b5b13
01fbdb93
02010513
02c10713
00072783
ffc72603
ffc70713
00379793
01d65613
00c7e7b3
00f72223
fee512e3
02012483
000087b7
fff78793
00349493
02912023
02fb1063
02812603
02412783
00c7e7b3
02c12603
00c7e7b3
0097e7b3
00079463
001bcb93
416405b3
113b94e3
2eb05463
01412c03
01812b83
01c12a83
0a0b1a63
02412603
02812783
02c12803
00f666b3
0106e6b3
0096e6b3
00069e63
03212823
03812a23
03712c23
03512e23
00058413
2ec0006f
fff58693
04069863
009904b3
01860633
02912823
0124b4b3
00960733
02e12a23
01863633
00973733
00e66633
017787b3
00c78733
02e12c23
0177b7b3
00c73733
00e7e7b3
01580833
010787b3
00100413
19c0006f
000087b7
fff78793
f8f586e3
07400793
04d7da63
02012623
02012423
02012223
00100793
11c0006f
000087b7
fff78793
00f41c63
03212823
03812a23
03712c23
03512e23
2500006f
02c12783
000806b7
00d7e7b3
02f12623
07400793
fab7cce3
00058693
4056d793
00070593
00000493
00000613
02f61e63
01f6f693
00279593
04069263
00300613
40f60633
00b70833
00082803
00168693
00470713
ff072e23
fed656e3
00400713
40f707b3
06c0006f
0005a803
00160613
00458593
0104e4b3
fb5ff06f
04058613
00260633
fe062603
02000893
40d888b3
01161633
00c4e4b3
00300613
00b505b3
00000313
40f60633
00458593
12c34a63
00400713
00261613
40f707b3
04060713
00270633
02c12703
00d75733
fee62023
00400613
40f60633
00279793
00f50533
00261613
00000593
850e20ef
02012703
009037b3
00f767b3
02f12023
02012783
02412703
00f907b3
00ec0733
02f12823
0127b7b3
00f706b3
02d12a23
00f6b6b3
02812783
01873733
00d76733
00fb87b3
00e786b3
02d12c23
00e6b6b3
02c12703
0177b7b3
00d7e7b3
00ea8733
00e787b3
00080737
02f12e23
00e7f733
0e070863
fff80737
fff70713
00e7f7b3
02f12e23
03012783
00140413
03c10593
01f79713
03010793
0007a683
0047a603
00478793
0016d693
01f61613
00c6e6b3
fed7ae23
feb792e3
03c12783
0017d793
02f12e23
00e037b3
03012703
00f767b3
02f12823
000087b7
fff78793
08f41263
02012e23
02012c23
02012a23
02012823
0700006f
ffc5a803
0005ae03
00130313
00d85833
011e1e33
01c86833
01072023
00470713
ea9ff06f
02412a83
02812b83
02c12c03
40058063
408b0633
20041a63
01412703
01812783
01c12503
00f765b3
00a5e5b3
0125e5b3
18059063
02912823
03512a23
03712c23
03812e23
00060413
03012783
0077f713
04070463
00f7f713
00400693
02d70e63
03412703
00478793
02f12823
0047b793
00e78733
02e12a23
00f73733
03812783
00f707b3
02f12c23
00e7b7b3
03c12703
00e787b3
02f12e23
03c12783
00080737
00e7f733
02070463
00008737
00140413
fff70713
00e41463
0100106f
fff80737
fff70713
00e7f7b3
02f12e23
03010793
03c10613
0007a703
0047a683
00478793
00375713
01d69693
00d76733
fee7ae23
fef612e3
03c12703
000086b7
fff68793
00375713
02e12e23
02f41a63
03412603
03012783
00c7e7b3
03812603
00c7e7b3
00e7e7b3
00078c63
02d12e23
02012c23
02012a23
02012823
00000993
03c12783
01141413
01145413
00f11623
03012783
00f99993
0089e9b3
00fa2023
03412783
01311723
06c12083
00fa2223
03812783
06812403
06412483
00fa2423
00c12783
06012903
05c12983
00fa2623
05412a83
05012b03
04c12b83
04812c03
04412c83
000a0513
05812a03
07010113
00008067
fff60893
04089663
00990933
01570733
03212823
00993933
012706b3
02d12a23
01573733
0126b6b3
00d76733
017787b3
00e786b3
02d12c23
0177b7b3
00e6b6b3
00d7e7b3
01850533
00a787b3
bb1ff06f
000087b7
fff78793
e2f606e3
07400793
0517dc63
00012e23
00012c23
00012a23
00100793
1640006f
000087b7
fff78793
00fb1e63
02912823
03512a23
03712c23
03812e23
000b0413
e01ff06f
01c12783
00080737
00e7e7b3
00f12e23
07400793
fac7cae3
00060893
41f8d793
01f7f793
011787b3
4057d793
00068613
00000413
00000713
04f74663
00078593
0007d463
00000593
01f8f513
00279613
04051463
00300593
00000713
40f585b3
00c68533
00052503
00170713
00468693
fea6ae23
fee5d6e3
00400713
40f707b3
08c0006f
00062583
00170713
00460613
00b46433
fa5ff06f
80000737
01f70713
00e8f733
00075863
fff70713
fe076713
00170713
00259593
02000893
40e888b3
04058713
002705b3
fd05a703
00c80633
00000313
01171733
00e46433
00300713
40f70733
00460613
0ae34a63
00400693
40f687b3
01c12683
00271713
04070713
00270733
00a6d6b3
fcd72823
00400713
00000613
00f74663
40f70733
00271613
00279793
00f80533
00000593
bbde10ef
01012703
008037b3
00f767b3
00f12823
01012783
01412703
000b0413
00f487b3
00ea8733
02f12823
0097b7b3
00f706b3
02d12a23
00f6b6b3
01812783
01573733
00d76733
00fb87b3
00e786b3
02d12c23
00e6b6b3
01c12703
0177b7b3
00d7e7b3
00ec0733
00e787b3
b69ff06f
ffc62583
00062e03
00130313
00a5d5b3
011e1e33
01c5e5b3
00b6a023
00468693
f29ff06f
00008837
00140693
ffe80893
0116f8b3
01412503
01812583
01c12703
03010793
03c10613
14089863
00b566b3
00e6e6b3
0126e6b3
0a041863
00069c63
02912823
03512a23
03712c23
03812e23
bf1ff06f
017ae7b3
0187e7b3
0097e7b3
00079c63
03212823
02a12a23
02b12c23
02e12e23
bcdff06f
009904b3
01550ab3
02912823
0124b4b3
009a87b3
02f12a23
00aabab3
0097b7b3
00faeab3
01758bb3
015b87b3
02f12c23
00bbbbb3
0157b7b3
00fbebb3
01870733
00eb8bb3
000807b7
00fbf7b3
00079663
03712e23
b75ff06f
fff807b7
fff78793
00fbfbb3
03712e23
00100413
b5dff06f
00069e63
02912823
03512a23
03712c23
03812e23
fff80413
b41ff06f
017aeab3
018aeab3
009aeab3
000a9c63
03212823
02a12a23
02b12c23
02e12e23
fd9ff06f
03012e23
02012c23
02012a23
02012823
00060713
00072683
ffc72603
ffc70713
00369693
01d65613
00c6e6b3
00d72223
fee792e3
03012783
00008437
00000993
00379793
02f12823
fff40413
acdff06f
009904b3
01550ab3
02912823
0124b4b3
009a8833
03012a23
00aabab3
00983833
010aeab3
01758bb3
015b8533
02a12c23
00bbbbb3
01553533
00abebb3
01870733
00eb8bb3
03712e23
0007a703
0047a583
00478793
00175713
01f59593
00b76733
fee7ae23
fef612e3
00008737
fff70713
03c12783
00e68a63
0017d793
02f12e23
00068413
a45ff06f
02012e23
02012c23
02012a23
02012823
fe9ff06f
26b05863
01412c03
01812b83
01c12a83
0a0b1263
02412603
02812803
02c12783
010666b3
00f6e6b3
0096e6b3
f0068063
fff58893
04089c63
40990733
40cc06b3
00e935b3
00dc3533
40b686b3
00000593
00e97663
41860633
00163593
00a5e5b3
410b8633
00cbb533
40b60633
00058663
41780833
00183893
40fa87b3
00a8e5b3
40b787b3
00100413
1980006f
000087b7
fff78793
e8f58c63
07400793
0517d063
02012623
02012423
02012223
00100793
10c0006f
000087b7
fff78793
f0f40863
02c12783
000806b7
00d7e7b3
02f12623
07400793
fcb7c6e3
00058893
4058d793
00070613
00000493
00000693
04f69063
01f8f893
00279613
04089463
00300593
00000693
40f585b3
00c70833
00082803
00168693
00470713
ff072e23
fed5d6e3
00400713
40f707b3
06c0006f
00062583
00168693
00460613
00b4e4b3
fb1ff06f
04060693
002686b3
fe06a683
02000813
41180833
010696b3
00d4e4b3
00300693
00c50633
00000313
40f686b3
00460613
0cd34e63
00400713
00269693
40f707b3
04068713
002706b3
02c12703
01175733
fee6a023
00400613
40f60633
00279793
00f50533
00261613
00000593
f6ce10ef
02012703
009037b3
00f767b3
02f12023
02012703
02412603
40e90733
40cc06b3
00e937b3
00dc35b3
40f686b3
00000793
00e97663
41860633
00163793
02812503
00b7e7b3
00000593
40ab8633
00cbb833
40f60633
00078663
41750533
00153593
02c12783
0105e5b3
40fa87b3
40b787b3
02e12823
00080737
02d12a23
02f12e23
02c12c23
00e7f6b3
fe068a63
fff70713
00e7f7b3
02f12e23
5ac0006f
ffc62583
00062e03
00130313
0115d5b3
010e1e33
01c5e5b3
00b72023
00470713
f01ff06f
02412a83
02812c03
02c12c83
2c058063
408b0733
0a041a63
01412603
01812583
01c12783
00b66533
00f56533
01256533
02051063
02912823
03512a23
03812c23
03912e23
00070413
000b8993
f70ff06f
fff70893
04089c63
41248733
40ca86b3
00e4b533
00dab833
40a686b3
00000513
00e4f663
41560633
00163513
01056533
40bc0633
00cc3833
40a60633
00050663
418585b3
0015b893
40fc87b3
0108e5b3
40b787b3
000b8993
d6dff06f
000087b7
fff78793
f8f700e3
07400793
1f17ce63
00088713
0400006f
000087b7
fff78793
00fb1e63
02912823
03512a23
03812c23
03912e23
000b0413
f61ff06f
01c12783
00080637
00c7e7b3
00f12e23
07400793
1ae7cc63
41f75793
01f7f793
00e787b3
4057d793
00068593
00000413
00000613
04f64663
00078593
0007d463
00000593
01f77893
00279613
04089463
00300593
00000713
40f585b3
00c68533
00052503
00170713
00468693
fea6ae23
fee5d6e3
00400713
40f707b3
08c0006f
0005a503
00160613
00458593
00a46433
fa5ff06f
80000537
01f50513
00a77733
00075863
fff70713
fe076713
00170713
00259593
02000513
40e50533
04058713
002705b3
fd05a703
00c80633
00000313
00a71733
00e46433
00300713
40f70733
00460613
0ce34263
00400693
40f687b3
01c12683
00271713
04070713
00270733
0116d6b3
fcd72823
00400713
00000613
00f74663
40f70733
00271613
00279793
00f80533
00000593
c94e10ef
01012703
008037b3
00f767b3
00f12823
01012703
01412603
40e48733
40ca86b3
00e4b7b3
00dab5b3
40f686b3
00000793
00e4f663
41560633
00163793
01812503
00b7e7b3
00000593
40ac0633
00cc3833
40f60633
00078663
41850533
00153593
01c12783
0105e5b3
000b0413
40fc87b3
40b787b3
000b8993
d21ff06f
ffc62583
00062e03
00130313
0115d5b3
00ae1e33
01c5e5b3
00b6a023
00468693
f19ff06f
00012e23
00012c23
00012a23
00100793
f5dff06f
00008537
ffe50713
00140793
00e7f7b3
01812683
01412703
01c12603
1e079063
018ae7b3
00d765b3
0197e7b3
00c5e5b3
0097e7b3
0125e5b3
10041a63
02059463
02912823
03512a23
03812c23
03912e23
000b8993
c8079e63
00000413
00000993
c90ff06f
00079c63
03212823
02e12a23
02d12c23
02c12e23
c78ff06f
409907b3
41570333
00f93533
00673833
40a30533
00000593
00f97463
00133593
0105e5b3
41868833
0106beb3
40b80e33
00000893
00058463
00183893
01d8e8b3
419605b3
411585b3
000808b7
02b12e23
03c12c23
02a12a23
02f12823
0115f8b3
06088063
41248933
40ea8733
0124b7b3
00eabab3
40f70733
00000793
0124f463
00133793
0157eab3
40dc06b3
00dc3c33
00000793
415686b3
000a8463
00183793
40cc8633
0187e7b3
40f60633
02c12e23
02d12c23
02e12a23
03212823
c45ff06f
00a7e7b3
01c7e7b3
00b7e7b3
f0dff06f
03010813
04059e63
02079e63
02a12e23
02012c23
02012a23
02012823
03c10793
0007a703
ffc7a683
ffc78793
00371713
01d6d693
00d76733
00e7a223
fef812e3
881ff06f
02912823
03512a23
03812c23
03912e23
000b8993
fff50413
b48ff06f
00079c63
03212823
02e12a23
02d12c23
02c12e23
fe5ff06f
02a12e23
02012c23
02012a23
02012823
03c10793
0007a703
ffc7a683
ffc78793
00371713
01d6d693
00d76733
00e7a223
fef812e3
815ff06f
409907b3
41570e33
00f93833
01c738b3
410e0833
00000513
00f97463
001e3513
01156533
418688b3
0116bf33
40a88eb3
00000313
00050463
0018b313
01e36333
41960533
40650533
00080337
02a12e23
03d12c23
03012a23
02f12823
00657333
16030663
41248933
40ea8733
0124b7b3
00eabab3
40f70733
00000793
0124f463
001e3793
40dc06b3
0157eab3
00dc3c33
415686b3
000a8463
0018b593
40cc8633
0185e7b3
40f60633
02c12e23
02d12c23
02e12a23
03212823
000b8993
03c12503
12050063
5f1000ef
ff450493
41f4d793
01f7f793
009787b3
4057d793
01f4f593
40f006b3
12058a63
80000737
01f70713
00e4f733
00075863
fff70713
fe076713
00170713
00269693
02000513
40e50533
03010893
00c68713
00e88733
40d006b3
12e89263
03012703
fff78613
00279793
04078793
002787b3
00b71733
fee7a823
00160613
00261613
00000593
03010513
890e10ef
2084c263
408487b3
00178793
41f7d513
01f57513
00f50533
03010613
40555513
00060693
00000413
00000713
0ea74463
00050693
00055463
00000693
01f7f813
00251713
0e081263
00300693
00000793
40a686b3
00e605b3
0005a583
00178793
00460613
feb62e23
fef6d6e3
00400793
40a78533
12c0006f
0107e7b3
01d7e7b3
00a7e7b3
c80782e3
ee1ff06f
03812503
00050863
4cd000ef
02050513
ed9ff06f
03412503
00050863
4b9000ef
04050513
ec5ff06f
03012503
4a9000ef
06050513
eb5ff06f
03c10713
00269693
00300613
00d705b3
0005a583
fff60613
ffc70713
00b72223
fef656e3
fff78613
f01ff06f
00072603
ffc72803
00d70333
00b61633
00a85833
01066633
00c32023
ffc70713
ebdff06f
0006a583
00170713
00468693
00b46433
f09ff06f
800005b7
01f58593
00b7f7b3
0007d863
fff78793
fe07e793
00178793
00269693
02000593
40f585b3
04068793
002786b3
ff06a783
00000893
00b797b3
00f46433
03010793
00e78733
00300793
40a787b3
00470713
06f8c263
00400713
40a70533
03c12703
00279793
04078793
002787b3
01075733
fee7a823
00400793
00000613
00a7c663
40a787b3
00279613
03010793
00251513
00a78533
00000593
ec9e00ef
03012703
008037b3
00000413
00f767b3
02f12823
fc5fe06f
ffc72683
00072303
00188893
0106d6b3
00b31333
0066e6b3
00d62023
00460613
f79ff06f
03c12783
fff80737
fff70713
00e7f7b3
40940433
02f12e23
f85fe06f
02012e23
02012c23
02012a23
02012823
ff5fe06f
00052683
00852783
00c52703
00452603
fe010113
00d12023
00f12423
00d12823
00f12c23
00171693
000047b7
00c12223
00e12623
0116d693
ffe78613
00000513
00d65e63
01d78613
01f75893
00d65c63
80000537
fff54513
00a88533
02010113
00008067
01071713
01075713
00010637
06f78793
40d787b3
00c76733
4057d693
00e12e23
01f7f793
04078863
ffe68813
02000513
00269693
40f50533
02068693
00a71533
00000313
00000613
00183813
002686b3
05064463
00030463
00b12823
00261613
02060693
00268633
00f75733
fee62823
0180006f
00269693
02068793
002786b3
ff06a783
00f12823
01012503
f60886e3
40a00533
f65ff06f
ff06a583
00100313
00100613
00f5d5b3
00a5e5b3
fa5ff06f
fc010113
02912a23
02112e23
02812c23
03212823
03312623
00050493
12058063
41f5d793
00b7c433
40f40433
00040513
01f5d913
1e5000ef
05150793
000049b7
01e98993
4057d713
00812823
00012a23
00012c23
00012e23
01f7f793
40a989b3
02078c63
00200693
0cd71663
02000693
40f686b3
00d456b3
00d12e23
fff70613
00271713
02070713
00270733
00f41433
fe872823
0340006f
00300793
40e787b3
00279793
02078793
002787b3
ff07a783
00200613
00f12e23
00200793
00f71663
00812c23
00100613
00160613
00000593
00261613
01010513
c6de00ef
00090593
01c12783
00f59413
01346433
00f11623
01012783
00811723
03c12083
00f4a023
01412783
03812403
03012903
00f4a223
01812783
02c12983
00048513
00f4a423
00c12783
00f4a623
03412483
04010113
00008067
00300713
f45ff06f
00012e23
00012c23
00012a23
00012823
00000993
f91ff06f
00800737
fff70713
01755693
00a77633
01f55793
0ff6f693
0175d513
0ff00813
00b77733
0ff57513
01f5d593
01069863
06060c63
00200513
00008067
01051463
fe071ae3
06069463
00051463
04070a63
00060e63
00b79463
02d55263
00100513
02078e63
fff00513
00008067
fff00513
02058663
00058513
00008067
00a6da63
fff00513
00078c63
00078513
00008067
fcc766e3
00000513
fee664e3
00008067
fe060ee3
fb9ff06f
f8d50ce3
fa0514e3
fa0706e3
fa1ff06f
008007b7
fff78793
00a7f733
01755513
00b7f7b3
0ff57513
0175d593
0ff00693
0ff5f593
00d51663
00100513
00071a63
0ff00713
00000513
00e59463
00f03533
00008067
01465793
00c61713
7ff7f793
fc010113
00c75713
00178693
02812c23
02912a23
03212823
02112e23
03312623
00b12823
00e12a23
00012e23
00012c23
7fe6f693
00050913
00058413
01f65493
08068463
000046b7
c0068693
00d787b3
00475693
00d12e23
01c71713
0045d693
00d76733
01c59413
00e12c23
00812a23
00012823
00f49493
00f4e4b3
01012783
01c12703
00911723
00f92023
01412783
00e11623
03c12083
00f92223
01812783
03812403
03412483
00f92423
00c12783
02c12983
00090513
00f92623
03012903
04010113
00008067
00b76533
0e079263
fa0502e3
06070063
00070513
6e0000ef
00050993
03198713
40575793
01f77713
40f006b3
04070663
00269693
00c68613
02000513
01010893
40e50533
00c88633
40d006b3
06c89c63
fff78613
00279793
02078793
002787b3
00e41733
fee7a823
0380006f
688000ef
02050993
fa9ff06f
01c10713
00269693
00300613
00d705b3
0005a583
fff60613
ffc70713
00b72223
fef656e3
fff78613
00160613
00261613
00000593
01010513
971e00ef
000047b7
c0c78793
413787b3
eedff06f
00062583
ffc62803
00d60333
00e595b3
00a85833
0105e5b3
00b32023
ffc60613
f69ff06f
000087b7
02050863
01c71793
0045d693
00d7e7b3
00f12c23
00475713
000087b7
01c59413
00f76733
00812a23
00012823
00e12e23
fff78793
e8dff06f
0145d613
7ff67613
00c59793
00160713
0097d793
01d55693
7fe77713
00f6e6b3
01f5d593
00351793
0a070663
c8060713
0fe00813
0ce84263
08e04063
fe900513
12a74063
00800537
00a6e6b3
01e00513
40e50533
01f00813
02a84863
c8260613
00a7d533
00c797b3
00f037b3
00c696b3
00d7e7b3
00f567b3
00000713
0077f693
08068063
0e40006f
ffe00813
40e80833
02000893
0106d833
00000713
01150663
ca260613
00c69733
00f76733
00e03733
00e867b3
fc5ff06f
00651513
00a03533
00369693
01d7d793
00d566b3
00f6e7b3
fadff06f
00f6e7b3
00061663
00f037b3
f99ff06f
0ff00713
00078c63
00369693
020007b7
fd9ff06f
00000793
0ff00713
040006b7
00d7f6b3
00068e63
00170713
0ff00693
06d70463
fc0006b7
fff68693
00d7f7b3
0ff00693
0037d793
00d71863
00078663
004007b7
00000593
7f8006b7
01771713
00979793
00d77733
0097d793
00f76733
01f59513
00a76533
00008067
00100793
00000713
00f7f693
00400613
f8c688e3
00478793
f89ff06f
00000793
fa5ff06f
fd010113
00852783
02912223
00c52483
00052683
00452703
00f12423
00f12c23
01049793
0107d793
00d12023
00d12823
00149693
00912623
00f12e23
02112623
02812423
00e12223
00e12a23
0116d693
01f4d493
01010513
01c10793
0007a703
ffc7a603
ffc78793
00371713
01d65613
00c76733
00e7a223
fef512e3
01012583
00008637
00168713
00359593
ffe60613
00b12823
00c77733
1a070663
ffffc737
40070713
00e686b3
7fe00713
1ed74863
06d05463
01812603
01c12783
01412703
01c65513
00479793
00a7e7b3
00f12a23
00471793
00b7e7b3
01c75713
00461613
00f037b3
00c76733
00e7e7b3
01412703
0077f613
1a060a63
00f7f613
00400593
1ab60463
00478613
00f637b3
00f70733
00060793
1940006f
fcc00713
00e6da63
00012a23
00100793
00000693
fc1ff06f
01c12703
00080837
00050593
00e86833
03d00713
40d706b3
01012e23
4056d713
00000613
00000413
0005a883
00160613
00458593
01146433
fec718e3
01f6f693
00271593
02069863
00300613
40e60633
00b78833
00082803
00168693
00478793
ff07ae23
fed656e3
00400793
40e78733
0540006f
02058613
00260633
ff062603
02000313
40d30333
00661633
00c46433
00300613
00b505b3
00000e13
40e60633
00458593
04ce4663
00400793
00261613
40e78733
02060793
00278633
00d85833
ff062823
00400613
40e60633
00271713
00e50533
00261613
00000593
d6ce00ef
01012703
008037b3
00e7e7b3
f0dff06f
ffc5a883
0005ae83
001e0e13
00d8d8b3
006e9eb3
01d8e8b3
0117a023
00478793
f91ff06f
01412603
01812703
01c12503
00c767b3
00a7e7b3
00b7e7b3
00069863
00f037b3
00000713
e89ff06f
0c078663
00471793
01c65613
01c75713
00451513
004006b7
00f66633
00a76733
00d76733
ff867793
7ff00693
e59ff06f
00000713
00000793
7ff00693
00800637
00c77633
00060e63
00168693
7ff00613
08c68263
ff800637
fff60613
00c77733
01d71613
0037d793
00f667b3
7ff00613
00375713
00c69e63
00e7e7b3
00000713
00078863
00080737
00000793
00000493
01469693
7ff00637
00c71713
02c12083
02812403
00c75713
00c6f6b3
01f49493
00e6e6b3
0096e733
00078513
02412483
00070593
03010113
00008067
00000713
f69ff06f
00000713
00000793
f85ff06f
00050313
ff010113
00060513
00068893
00112623
00030613
00050693
00000713
00000793
00000813
0016fe13
00171e93
000e0c63
01060e33
010e3833
00e787b3
00f807b3
000e0813
01f65713
0016d693
00eee733
00161613
fc0698e3
00058663
dbdde0ef
00a787b3
00088a63
00030513
00088593
da9de0ef
00f507b3
00c12083
00080513
00078593
01010113
00008067
02060063
02000793
40c787b3
00f04c63
fe060613
00c5d533
00000713
00070593
00008067
00c5d733
00c55533
00f595b3
00b56533
fe9ff06f
02060063
02000793
40c787b3
00f04c63
fe060613
00c515b3
00000713
00070513
00008067
00c51733
00c595b3
00f55533
00a5e5b3
fe9ff06f
000107b7
02f57a63
10053793
0017c793
00379793
00025737
02000693
40f686b3
00f55533
c0870793
00a787b3
0007c503
40a68533
00008067
01000737
01000793
fce56ae3
01800793
fcdff06f
f7010113
08112623
08812423
08912223
09212023
07312e23
07412c23
07512a23
07612823
07712623
07812423
07912223
07a12023
05b12e23
200007b7
fff00713
000104b7
30e7a423
fff48493
3097a623
00600713
30e7a223
03e00513
c00e00ef
04001db7
9e4da783
00025d37
04000bb7
0087a503
00000413
00000993
824df0ef
e3cd0793
00f12423
ffffe7b7
bfe78793
000b8b93
04259937
07f00a13
00800b13
03f00c13
00a00c93
02000a93
00f12623
af9de0ef
02051a63
b3d94783
00078463
cd5dd0ef
cd8de0ef
009477b3
00140413
fe0790e3
41045793
20000737
00f72823
ac9de0ef
fc050ae3
af1de0ef
00050793
03450a63
03650863
053c4063
05950463
00d00713
04e50063
04098713
01010693
00d70733
fca70023
00198993
afdde0ef
f99ff06f
f8098ae3
00078513
fff98993
ae9de0ef
f85ff06f
00700513
addde0ef
f79ff06f
04098793
01010713
00e789b3
00a00513
fc098023
ac1de0ef
01014783
01010d13
01579863
001d4703
001d0d13
ff570ce3
02000593
000d0513
ff8e00ef
00812983
00050663
00050023
00150993
004ba583
000d0513
91de00ef
06050863
00cba583
000d0513
90de00ef
04050e63
014ba583
000d0513
8fde00ef
06050e63
01cba583
000d0513
8ede00ef
06050a63
000d4703
00d00693
04e6f663
000257b7
000d0593
e0478513
a1ce00ef
03e00513
a6ce00ef
9e4da783
00000993
0087a503
ea1de0ef
eb5ff06f
00100513
00351793
00fb87b3
0007a783
00098513
000780e7
fcdff06f
00c12783
40e7d733
00177713
fa070ee3
fa9ff06f
00200513
fd1ff06f
00300513
fc9ff06f
00000793
00078863
00009537
d5450513
92cf406f
00008067
00000190
00024e6c
00000458
00024e74
00000d88
00024e7c
00000168
00024e84
00000000
0400030c
04000374
040003dc
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000001
00000000
abcd330e
e66d1234
0005deec
0000000b
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
04000448
04000448
04000450
04000450
04000458
04000458
04000460
04000460
04000468
04000468
04000470
04000470
04000478
04000478
04000480
04000480
04000488
04000488
04000490
04000490
04000498
04000498
040004a0
040004a0
040004a8
040004a8
040004b0
040004b0
040004b8
040004b8
040004c0
040004c0
040004c8
040004c8
040004d0
040004d0
040004d8
040004d8
040004e0
040004e0
040004e8
040004e8
040004f0
040004f0
040004f8
040004f8
04000500
04000500
04000508
04000508
04000510
04000510
04000518
04000518
04000520
04000520
04000528
04000528
04000530
04000530
04000538
04000538
04000540
04000540
04000548
04000548
04000550
04000550
04000558
04000558
04000560
04000560
04000568
04000568
04000570
04000570
04000578
04000578
04000580
04000580
04000588
04000588
04000590
04000590
04000598
04000598
040005a0
040005a0
040005a8
040005a8
040005b0
040005b0
040005b8
040005b8
040005c0
040005c0
040005c8
040005c8
040005d0
040005d0
040005d8
040005d8
040005e0
040005e0
040005e8
040005e8
040005f0
040005f0
040005f8
040005f8
04000600
04000600
04000608
04000608
04000610
04000610
04000618
04000618
04000620
04000620
04000628
04000628
04000630
04000630
04000638
04000638
04000640
04000640
04000648
04000648
04000650
04000650
04000658
04000658
04000660
04000660
04000668
04000668
04000670
04000670
04000678
04000678
04000680
04000680
04000688
04000688
04000690
04000690
04000698
04000698
040006a0
040006a0
040006a8
040006a8
040006b0
040006b0
040006b8
040006b8
040006c0
040006c0
040006c8
040006c8
040006d0
040006d0
040006d8
040006d8
040006e0
040006e0
040006e8
040006e8
040006f0
040006f0
040006f8
040006f8
04000700
04000700
04000708
04000708
04000710
04000710
04000718
04000718
04000720
04000720
04000728
04000728
04000730
04000730
04000738
04000738
04000740
04000740
04000748
04000748
04000750
04000750
04000758
04000758
04000760
04000760
04000768
04000768
04000770
04000770
04000778
04000778
04000780
04000780
04000788
04000788
04000790
04000790
04000798
04000798
040007a0
040007a0
040007a8
040007a8
040007b0
040007b0
040007b8
040007b8
040007c0
040007c0
040007c8
040007c8
040007d0
040007d0
040007d8
040007d8
040007e0
040007e0
040007e8
040007e8
040007f0
040007f0
040007f8
040007f8
04000800
04000800
04000808
04000808
04000810
04000810
04000818
04000818
04000820
04000820
04000828
04000828
04000830
04000830
04000838
04000838
04000840
04000840
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
000166e8
0000c314
00000000
00023c00
00024f74
00024e3c
00024e3c
00024e3c
00024e3c
00024e3c
00024e3c
00024e3c
00024e3c
00024e3c
ffffffff
ffffffff
ffffffff
0000ffff
53410001
00494943
00000000
00000000
00000000
00000000
00000000
00000000
53410000
00494943
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000040
ffffbfc3
00003fc0
00000001
00000000
00000000
00000001
ffffffff
ffffffff
00000101
04000020
ffffffff
00020000
000000ff
00000010
00000000
00527a03
01017c01
00020d1b
00000048
00000018
fc01b1bc
000005c0
300e4400
8105936c
89028801
94049203
96079506
98099708
030b990a
c10a0254
c944c844
d444d344
d644d544
d844d744
d24cd944
44000e44
0000000b
0000004c
00000064
fc01b730
000004d0
300e4400
89028870
92018103
94059304
96079506
98099708
9a0b990a
010c030c
c844c10a
d244c944
d444d344
d644d544
d844d744
da44d944
44000e44
0000000b
00000000
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
000005cc
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000784
0000078c
00000738
00000730
00000728
00000720
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000700
00000784
0000078c
00000738
00000730
00000728
00000720
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005ec
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
00000764
00000758
0000074c
00000740
00000714
00000708
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
000005f8
00000764
00000758
0000074c
00000740
00000714
00000708
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007cc
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
00000800
00000808
000007e0
000007f0
000007f8
000007e8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
000007d8
00000800
00000808
000007e0
000007f0
000007f8
000007e8
b0a4f9c0
f8829299
83889080
8e86a1c6
00003308
00003504
00003504
00003504
00003504
00003b28
00003504
00003504
00003504
00003504
00003504
00003520
00003520
00003520
00003520
00003520
00003520
00003520
00003520
00003520
00003520
00003504
00003504
00003504
00003504
00003504
00003504
00003504
00003548
00003504
00003990
000039dc
00003548
00003548
00003548
00003504
00003504
00003504
00003504
000038b0
00003504
00003504
000039b4
00003504
00003504
00003504
000039a4
00003504
00003504
00003504
00003504
000038d4
00003504
00003504
00003a34
00003504
00003504
00003504
00003504
00003504
00003548
00003504
00003994
000039e0
00003548
00003548
00003548
00003a04
00003a54
000038b0
00003504
00003a88
00003aa8
00003ad8
000039b8
00003b20
00003504
00003504
000039a8
000038c8
00003a24
00003504
00003504
000038d4
00003504
000038c8
000040d4
0000401c
000040d4
0000401c
0000401c
00004358
000040ac
000040ac
000040ac
000040ac
000040ac
000040ac
000040ac
000040ac
000040ac
0000401c
0000401c
0000401c
0000401c
0000401c
0000401c
0000401c
000040c4
0000401c
0000401c
0000401c
000042d4
000042c4
0000401c
0000401c
00004118
0000401c
0000401c
0000401c
0000401c
000040e4
0000401c
0000401c
0000401c
0000401c
0000401c
00004348
0000401c
0000401c
0000401c
0000401c
00004338
0000401c
0000401c
0000401c
0000401c
0000401c
0000401c
0000401c
000040c4
0000401c
0000401c
0000401c
000042d4
000042c4
0000401c
0000401c
00004118
0000401c
0000401c
0000401c
0000401c
000040e4
0000401c
0000401c
0000401c
0000401c
0000401c
00004348
0000401c
0000401c
0000401c
0000401c
00004338
000045ac
000044a0
000045ac
000044a0
000044a0
000045d4
0000457c
0000457c
0000457c
0000457c
0000457c
0000457c
0000457c
000045bc
000045bc
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
0000446c
0000446c
0000446c
0000446c
0000446c
0000446c
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
00004590
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
0000446c
0000446c
0000446c
0000446c
0000446c
0000446c
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
000044a0
00004590
0001000a
00030002
00050004
00070006
00090008
000b000a
000d000c
000f000e
00000010
000067dc
00006018
00006018
000067d0
00006018
00006018
00006018
00006204
00006018
00006018
00006648
00006770
00006018
00006660
0000678c
00006018
00006780
00005fe8
00005fe8
00005fe8
00005fe8
00005fe8
00005fe8
00005fe8
00005fe8
00005fe8
00006018
00006018
00006018
00006018
00006018
00006018
00006018
0000627c
00006018
000065a0
0000686c
0000627c
0000627c
0000627c
00006018
00006018
00006018
00006018
00006860
00006018
00006018
000067f4
00006018
00006018
00006018
000065c8
00006018
0000682c
00006018
00006018
0000723c
00006018
00006018
00006018
00006018
00006018
00006018
00006018
00006018
0000627c
00006018
000065a0
000070fc
0000627c
0000627c
0000627c
0000675c
000070fc
00006244
00006018
000066b4
00006018
0000666c
00007250
000066c8
00006244
00006018
000065c8
0000623c
000071d0
00006018
00006018
000071dc
00006018
0000623c
00008044
0000796c
0000796c
0000796c
0000802c
00008038
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000796c
0000802c
00008038
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
20202000
20202020
28282020
20282828
20202020
20202020
20202020
20202020
10108820
10101010
10101010
10101010
04040410
04040404
10040404
10101010
41411010
41414141
01010101
01010101
01010101
01010101
01010101
10101010
42421010
42424242
02020202
02020202
02020202
02020202
02020202
10101010
00000020
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
3fff8000
4a926576
153f804a
979ac94c
52028a20
7525c460
ce526a32
28ce329a
5de4a74d
3b5dc53d
5a929e8b
50ce526c
3d28f18b
0c17650d
75868175
4d48c976
58f89c66
5c54bc50
91c6cc65
a0aea60e
46a3e319
eab7851e
901b98fe
de8dddbb
ebfb9df9
4351aa7e
01370235
336c36b1
8cdfc66f
47c980e9
41a893ba
25fb50f8
6b71c76b
a6d53cbf
1f49ffcf
40d3c278
00000000
00000000
b59df020
ada82b70
40699dc5
00000000
00000000
00000000
c9bf0400
40348e1b
00000000
00000000
00000000
20000000
4019bebc
00000000
00000000
00000000
00000000
400c9c40
00000000
00000000
00000000
00000000
4005c800
00000000
00000000
00000000
00000000
4002a000
cffc2030
8123a1c3
9fde2de3
04c8d2ce
0ad8a6dd
d2cb8264
12d4f2ea
2de44925
534f3436
256bceae
f698f53f
01586bd3
c0bd87a6
82a5da57
32b5a2a6
04d4e731
d332e3f2
d21c7132
ee32db23
395a9049
5308a23e
1155fefb
1939fa91
4325637a
3cacc031
dbdee26d
b3f6d05d
e4a0ac7c
467c64bc
3e55ddd0
62242a20
98d747b3
e9a53f23
ea27a539
3f2aa87f
4af20b5b
18eda581
94ba67de
1ead4539
3f94cfb1
a9b3bf71
be687989
e15b4c2e
94bec44d
3fc9e695
7c3d3d4d
0d2b36ba
cefcfdc2
77118461
3fe4abcc
a4a8c155
6113404e
652bd3c3
1758e219
3ff1d1b7
70a3d70a
a3d70a3d
d70a3d70
0a3d70a3
3ff8a3d7
cccccccd
cccccccc
cccccccc
cccccccc
3ffbcccc
fffeffff
fff8fffc
ffe0fff0
ff80ffc0
fe00ff00
f800fc00
e000f000
8000c000
00000000
00000005
00000019
0000007d
00000000
00000000
3ff00000
00000000
40240000
00000000
40590000
00000000
408f4000
00000000
40c38800
00000000
40f86a00
00000000
412e8480
00000000
416312d0
00000000
4197d784
00000000
41cdcd65
20000000
4202a05f
e8000000
42374876
a2000000
426d1a94
e5400000
42a2309c
1e900000
42d6bcc4
26340000
430c6bf5
37e08000
4341c379
85d8a000
43763457
674ec800
43abc16d
60913d00
43e158e4
78b58c40
4415af1d
d6e2ef50
444b1ae4
064dd592
4480f0cf
c7e14af6
44b52d02
79d99db4
44ea7843
97d889bc
3c9cd2b2
d5a8a733
3949f623
44f4a73d
32a50ffd
cf8c979d
255bba08
64ac6f43
0ac80628
37e08000
4341c379
b5056e17
4693b8b5
e93ff9f5
4d384f03
f9301d32
5a827748
7f73bf3c
75154fdd
0000e618
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e66c
0000e66c
0000e66c
0000e66c
0000e66c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e66c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000e53c
0000f2bc
0000e53c
0000e600
0000f570
0000f550
0000f5a0
0000f598
0000f588
0000f550
00000035
fffffbce
000003cb
00000001
00000000
00000034
fffffbce
000003cb
00000001
00000000
97d889bc
3c9cd2b2
d5a8a733
3949f623
44f4a73d
32a50ffd
cf8c979d
255bba08
64ac6f43
11680628
00010420
000103cc
00010488
00010460
00010440
000103cc
00010420
00010f38
000110a8
000110a8
000110a8
000110a8
00011518
000110a8
000110a8
000110a8
000110a8
000110a8
000110b8
000110b8
000110b8
000110b8
000110b8
000110b8
000110b8
000110b8
000110b8
000110b8
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
00011478
00011454
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
000110ec
000110a8
000110a8
000112f0
000110a8
000110a8
000110a8
00011444
000110a8
000110a8
000110a8
000110a8
00011104
000110a8
000110a8
000113cc
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
000110a8
00012178
00012180
000110a8
000110a8
000110a8
00011408
00011428
000110ec
000110a8
000113e8
0001148c
000114b0
00012170
000114e0
000110a8
000110a8
000114ec
000110e0
000114f8
000110a8
000110a8
00011104
000110a8
000110e0
00011a94
000119f8
00011a94
000119f8
000119f8
00011ac0
00011a60
00011a60
00011a60
00011a60
00011a60
00011a60
00011a60
00011aa4
00011aa4
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119c4
000119c4
000119c4
000119c4
000119c4
000119c4
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
00011a78
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119c4
000119c4
000119c4
000119c4
000119c4
000119c4
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
000119f8
00011a78
0001000a
00030002
00050004
00070006
00090008
000b000a
000d000c
000f000e
00000010
000131c0
00012a2c
00012a2c
000131b4
00012a2c
00012a2c
00012a2c
00012bd0
00012a2c
00012a2c
0001300c
00013228
00012a2c
00013024
000131e4
00012a2c
000131d8
000129fc
000129fc
000129fc
000129fc
000129fc
000129fc
000129fc
000129fc
000129fc
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012c4c
00012a2c
00012fe4
00013238
00012c4c
00012c4c
00012c4c
00012a2c
00012a2c
00012a2c
00012a2c
000131a8
00012a2c
00012a2c
00013128
00012a2c
00012a2c
00012a2c
00012f64
00012a2c
00013174
00012a2c
00012a2c
00013c94
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012a2c
00012c4c
00012a2c
00012fe4
00013b2c
00012c4c
00012c4c
00012c4c
00013160
00013b2c
00012c14
00012a2c
00013080
00012a2c
00013030
00013ca8
00013094
00012c14
00012a2c
00012f64
00012c0c
00013be8
00012a2c
00012a2c
00013bf4
00012a2c
00012c0c
000146b0
000143f4
000143f4
000143f4
00014698
000146a4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
000143f4
00014698
000146a4
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
00015be0
00015634
00015634
00015bd4
00015634
00015634
00015634
000157f0
00015634
00015634
00015b4c
00015c44
00015634
00015b70
00015c04
00015634
00015bf8
000155fc
000155fc
000155fc
000155fc
000155fc
000155fc
000155fc
000155fc
000155fc
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015af8
00015840
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015938
00015634
00015634
00015634
00015ab8
00015634
00015ba4
00015634
00015634
000163f0
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015634
00015af8
00015844
00015634
00015634
00015634
00015b90
00015844
00015834
00015634
00015b7c
00015634
00015c8c
0001593c
00015c54
00015834
00015634
00015ab8
0001582c
0001638c
00015634
00015634
00016394
00015634
0001582c
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
13121110
17161514
00001918
00000000
1c1b1a00
001f1e1d
00000000
00000000
00000000
00000000
00000000
00000000
1c1b1a00
001f1e1d
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00024f74
00024e3c
040009f0
00018290
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000182ec
000182ec
000182ec
000182ec
000182ec
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000182ec
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
000181a4
00018ef0
000181a4
00018278
00000000
00000003
00000005
00000007
0000000a
0000000c
0000000e
00000011
00000013
00000015
00000018
0000001a
0000001c
0000001f
00000021
00000023
00000026
00000028
0000002a
0000002d
0000002f
00000031
00000034
0001a8e0
0001a2f0
0001a2f0
0001a8d4
0001a2f0
0001a2f0
0001a2f0
0001a45c
0001a2f0
0001a2f0
0001a8b4
0001a8a4
0001a2f0
0001a4c0
0001a864
0001a2f0
0001a6f8
0001a2b8
0001a2b8
0001a2b8
0001a2b8
0001a2b8
0001a2b8
0001a2b8
0001a2b8
0001a2b8
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a594
0001a790
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a75c
0001a2f0
0001a2f0
0001a2f0
0001a540
0001a2f0
0001a72c
0001a2f0
0001a2f0
0001afd4
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a2f0
0001a594
0001a5c0
0001a2f0
0001a2f0
0001a2f0
0001a718
0001a5c0
0001a4a4
0001a2f0
0001a704
0001a2f0
0001a6b8
0001b01c
0001a644
0001a4a4
0001a2f0
0001a540
0001a49c
0001af6c
0001a2f0
0001a2f0
0001af74
0001a2f0
0001a49c
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
0001d4fc
0001d5dc
0001d50c
0001d5dc
0001d5e8
0001d5dc
0001d50c
0001d4fc
0001d4fc
0001d5e8
0001d50c
0001d4d4
0001d4d4
0001d4d4
0001d514
02020100
03030303
04040404
04040404
05050505
05050505
05050505
05050505
06060606
06060606
06060606
06060606
06060606
06060606
06060606
06060606
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
3a6d756e
2c642520
6d617320
72656c70
3a657461
2c642520
74696220
25203a73
00000a64
0000002d
00006425
736d656d
203a7465
65726e75
6e676f63
64657a69
65706f20
646e6172
73252720
00000a27
64616552
20676e69
62206425
73657479
206f7420
626d656d
6b636f6c
0a642520
00000000
626d654d
6b636f6c
3a444920
20642520
2074756f
7220666f
65676e61
616d202c
73692078
0a642520
00000000
62616e55
7420656c
6c61206f
61636f6c
6d206574
726f6d65
6d202c79
6f6c6c61
20292863
75746572
64656e72
4c554e20
00000a4c
20202020
20202020
20202020
20202020
0000000d
65646956
6e69206f
61697469
657a696c
00000064
203a7325
6d6d6f63
20646e61
20746f6e
6e756f66
00000a64
79616c70
6e75203a
6f636572
7a696e67
6f206465
61726570
2720646e
0a277325
00000000
79616c50
203a676e
69647561
6f73206f
65637275
2c64253d
64697620
73206f65
6372756f
64253d65
0000000a
6f686365
00000000
736d656d
00007465
79616c70
00000000
706f7473
00000000
646c2565
00000000
00464e49
00666e69
004e414e
006e616e
33323130
37363534
62613938
66656463
00000000
33323130
37363534
42413938
46454443
00000000
6c756e28
0000296c
00000030
6e492d20
696e6966
00207974
666e4920
74696e69
00002079
004e614e
00642545
6c6c6142
7320636f
65636375
64656465
00000000
6d6f682f
62752f65
75746e75
636f442f
6e656d75
722f7374
76637369
756e672d
6f6f742d
6168636c
722f6e69
76637369
77656e2d
2f62696c
6c77656e
6c2f6269
2f636269
6c647473
6c2f6269
616f7464
0000632e
4e614e20
00000020
00000043
49534f50
00000058
0000002e
6d6f682f
62752f65
75746e75
636f442f
6e656d75
722f7374
76637369
756e672d
6f6f742d
6168636c
722f6e69
76637369
77656e2d
2f62696c
6c77656e
6c2f6269
2f636269
6c647473
6d2f6269
63657270
0000632e
0000666e
74696e69
00000079
00006e61
7566202c
6974636e
203a6e6f
00000000
65737361
6f697472
2522206e
66202273
656c6961
66203a64
20656c69
22732522
696c202c
2520656e
25732564
00000a73
6d6f682f
62752f65
75746e75
636f442f
6e656d75
722f7374
76637369
756e672d
6f6f742d
6168636c
722f6e69
76637369
77656e2d
2f62696c
6c77656e
6c2f6269
2f636269
6c647473
672f6269
616f7464
7465672d
2e786568
00000063
6d6f682f
62752f65
75746e75
636f442f
6e656d75
722f7374
76637369
756e672d
6f6f742d
6168636c
722f6e69
76637369
77656e2d
2f62696c
6c77656e
6c2f6269
2f636269
6c647473
732f6269
6f747274
632e6764
00000000
04000020
00000000
00000000
3ff00000
00000000
40240000
7fc00000
00000000
00000000
43500000
00000000
3fe00000
00000000
40000000
ffc00000
41dfffff
94a03595
3fdfffff
35afe535
3fe00000
94a03595
3fcfffff
00000000
39500000
ffffffff
7fefffff
7f7fffff
00000000
99999999
19999999
00000000
7ff80000
9ee75616
3cc203af
00000110
00022648
000000c8
