-- system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		av_dac_external_interface_acknowledge  : in    std_logic                     := '0';             --  av_dac_external_interface.acknowledge
		av_dac_external_interface_irq          : in    std_logic                     := '0';             --                           .irq
		av_dac_external_interface_address      : out   std_logic_vector(2 downto 0);                     --                           .address
		av_dac_external_interface_bus_enable   : out   std_logic;                                        --                           .bus_enable
		av_dac_external_interface_byte_enable  : out   std_logic_vector(3 downto 0);                     --                           .byte_enable
		av_dac_external_interface_rw           : out   std_logic;                                        --                           .rw
		av_dac_external_interface_write_data   : out   std_logic_vector(31 downto 0);                    --                           .write_data
		av_dac_external_interface_read_data    : in    std_logic_vector(31 downto 0) := (others => '0'); --                           .read_data
		av_uart_external_interface_acknowledge : in    std_logic                     := '0';             -- av_uart_external_interface.acknowledge
		av_uart_external_interface_irq         : in    std_logic                     := '0';             --                           .irq
		av_uart_external_interface_address     : out   std_logic_vector(2 downto 0);                     --                           .address
		av_uart_external_interface_bus_enable  : out   std_logic;                                        --                           .bus_enable
		av_uart_external_interface_byte_enable : out   std_logic_vector(3 downto 0);                     --                           .byte_enable
		av_uart_external_interface_rw          : out   std_logic;                                        --                           .rw
		av_uart_external_interface_write_data  : out   std_logic_vector(31 downto 0);                    --                           .write_data
		av_uart_external_interface_read_data   : in    std_logic_vector(31 downto 0) := (others => '0'); --                           .read_data
		av_vga_external_interface_acknowledge  : in    std_logic                     := '0';             --  av_vga_external_interface.acknowledge
		av_vga_external_interface_irq          : in    std_logic                     := '0';             --                           .irq
		av_vga_external_interface_address      : out   std_logic_vector(3 downto 0);                     --                           .address
		av_vga_external_interface_bus_enable   : out   std_logic;                                        --                           .bus_enable
		av_vga_external_interface_byte_enable  : out   std_logic_vector(3 downto 0);                     --                           .byte_enable
		av_vga_external_interface_rw           : out   std_logic;                                        --                           .rw
		av_vga_external_interface_write_data   : out   std_logic_vector(31 downto 0);                    --                           .write_data
		av_vga_external_interface_read_data    : in    std_logic_vector(31 downto 0) := (others => '0'); --                           .read_data
		clk_clk                                : in    std_logic                     := '0';             --                        clk.clk
		clk_sdram_clk                          : out   std_logic;                                        --                  clk_sdram.clk
		disp0_export                           : out   std_logic_vector(7 downto 0);                     --                      disp0.export
		disp1_export                           : out   std_logic_vector(7 downto 0);                     --                      disp1.export
		disp2_export                           : out   std_logic_vector(7 downto 0);                     --                      disp2.export
		disp3_export                           : out   std_logic_vector(7 downto 0);                     --                      disp3.export
		disp4_export                           : out   std_logic_vector(7 downto 0);                     --                      disp4.export
		disp5_export                           : out   std_logic_vector(7 downto 0);                     --                      disp5.export
		leds_export                            : out   std_logic_vector(9 downto 0);                     --                       leds.export
		rst_reset_n                            : in    std_logic                     := '0';             --                        rst.reset_n
		sdram_addr                             : out   std_logic_vector(12 downto 0);                    --                      sdram.addr
		sdram_ba                               : out   std_logic_vector(1 downto 0);                     --                           .ba
		sdram_cas_n                            : out   std_logic;                                        --                           .cas_n
		sdram_cke                              : out   std_logic;                                        --                           .cke
		sdram_cs_n                             : out   std_logic;                                        --                           .cs_n
		sdram_dq                               : inout std_logic_vector(15 downto 0) := (others => '0'); --                           .dq
		sdram_dqm                              : out   std_logic_vector(1 downto 0);                     --                           .dqm
		sdram_ras_n                            : out   std_logic;                                        --                           .ras_n
		sdram_we_n                             : out   std_logic;                                        --                           .we_n
		sys_clk                                : out   std_logic                                         --                        sys.clk
	);
end entity system;

architecture rtl of system is
	component system_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component system_altpll_0;

	component system_av_dac is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			avalon_address     : in  std_logic                     := 'X';             -- address
			avalon_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avalon_chipselect  : in  std_logic                     := 'X';             -- chipselect
			avalon_read        : in  std_logic                     := 'X';             -- read
			avalon_write       : in  std_logic                     := 'X';             -- write
			avalon_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_waitrequest : out std_logic;                                        -- waitrequest
			avalon_irq         : out std_logic;                                        -- irq
			acknowledge        : in  std_logic                     := 'X';             -- export
			irq                : in  std_logic                     := 'X';             -- export
			address            : out std_logic_vector(2 downto 0);                     -- export
			bus_enable         : out std_logic;                                        -- export
			byte_enable        : out std_logic_vector(3 downto 0);                     -- export
			rw                 : out std_logic;                                        -- export
			write_data         : out std_logic_vector(31 downto 0);                    -- export
			read_data          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component system_av_dac;

	component system_av_vga is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			avalon_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avalon_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avalon_chipselect  : in  std_logic                     := 'X';             -- chipselect
			avalon_read        : in  std_logic                     := 'X';             -- read
			avalon_write       : in  std_logic                     := 'X';             -- write
			avalon_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_waitrequest : out std_logic;                                        -- waitrequest
			avalon_irq         : out std_logic;                                        -- irq
			acknowledge        : in  std_logic                     := 'X';             -- export
			irq                : in  std_logic                     := 'X';             -- export
			address            : out std_logic_vector(3 downto 0);                     -- export
			bus_enable         : out std_logic;                                        -- export
			byte_enable        : out std_logic_vector(3 downto 0);                     -- export
			rw                 : out std_logic;                                        -- export
			write_data         : out std_logic_vector(31 downto 0);                    -- export
			read_data          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component system_av_vga;

	component system_code_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_code_ram;

	component system_disp_7_seg is
		port (
			pio_disp_0_clk_clk                    : in  std_logic                     := 'X';             -- clk
			pio_disp_0_external_connection_export : out std_logic_vector(7 downto 0);                     -- export
			pio_disp_0_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			pio_disp_0_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pio_disp_0_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			pio_disp_0_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_disp_0_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			pio_disp_0_s1_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			pio_disp_1_clk_clk                    : in  std_logic                     := 'X';             -- clk
			pio_disp_1_external_connection_export : out std_logic_vector(7 downto 0);                     -- export
			pio_disp_1_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			pio_disp_1_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pio_disp_1_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			pio_disp_1_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_disp_1_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			pio_disp_1_s1_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			pio_disp_2_clk_clk                    : in  std_logic                     := 'X';             -- clk
			pio_disp_2_external_connection_export : out std_logic_vector(7 downto 0);                     -- export
			pio_disp_2_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			pio_disp_2_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pio_disp_2_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			pio_disp_2_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_disp_2_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			pio_disp_2_s1_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			pio_disp_3_clk_clk                    : in  std_logic                     := 'X';             -- clk
			pio_disp_3_external_connection_export : out std_logic_vector(7 downto 0);                     -- export
			pio_disp_3_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			pio_disp_3_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pio_disp_3_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			pio_disp_3_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_disp_3_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			pio_disp_3_s1_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			pio_disp_4_clk_clk                    : in  std_logic                     := 'X';             -- clk
			pio_disp_4_external_connection_export : out std_logic_vector(7 downto 0);                     -- export
			pio_disp_4_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			pio_disp_4_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pio_disp_4_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			pio_disp_4_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_disp_4_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			pio_disp_4_s1_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			pio_disp_5_clk_clk                    : in  std_logic                     := 'X';             -- clk
			pio_disp_5_external_connection_export : out std_logic_vector(7 downto 0);                     -- export
			pio_disp_5_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			pio_disp_5_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pio_disp_5_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			pio_disp_5_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pio_disp_5_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			pio_disp_5_s1_readdata                : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component system_disp_7_seg;

	component system_pio_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component system_pio_leds;

	component riscv_mk1 is
		port (
			o_av_addr        : out std_logic_vector(29 downto 0);                    -- address
			o_av_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			o_av_read        : out std_logic;                                        -- read
			o_av_write       : out std_logic;                                        -- write
			i_av_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			o_av_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			i_av_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_clk            : in  std_logic                     := 'X';             -- clk
			i_rst            : in  std_logic                     := 'X'              -- reset
		);
	end component riscv_mk1;

	component system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_sdram;

	component system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component system_timer_0;

	component system_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                               : in  std_logic                     := 'X';             -- clk
			riscv_mk1_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			riscv_mk1_0_avalon_master_address             : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			riscv_mk1_0_avalon_master_waitrequest         : out std_logic;                                        -- waitrequest
			riscv_mk1_0_avalon_master_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			riscv_mk1_0_avalon_master_read                : in  std_logic                     := 'X';             -- read
			riscv_mk1_0_avalon_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			riscv_mk1_0_avalon_master_write               : in  std_logic                     := 'X';             -- write
			riscv_mk1_0_avalon_master_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_dac_avalon_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			av_dac_avalon_slave_write                     : out std_logic;                                        -- write
			av_dac_avalon_slave_read                      : out std_logic;                                        -- read
			av_dac_avalon_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_dac_avalon_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			av_dac_avalon_slave_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			av_dac_avalon_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			av_dac_avalon_slave_chipselect                : out std_logic;                                        -- chipselect
			av_uart_avalon_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			av_uart_avalon_slave_write                    : out std_logic;                                        -- write
			av_uart_avalon_slave_read                     : out std_logic;                                        -- read
			av_uart_avalon_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_uart_avalon_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			av_uart_avalon_slave_byteenable               : out std_logic_vector(3 downto 0);                     -- byteenable
			av_uart_avalon_slave_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			av_uart_avalon_slave_chipselect               : out std_logic;                                        -- chipselect
			av_vga_avalon_slave_address                   : out std_logic_vector(1 downto 0);                     -- address
			av_vga_avalon_slave_write                     : out std_logic;                                        -- write
			av_vga_avalon_slave_read                      : out std_logic;                                        -- read
			av_vga_avalon_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_vga_avalon_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			av_vga_avalon_slave_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			av_vga_avalon_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			av_vga_avalon_slave_chipselect                : out std_logic;                                        -- chipselect
			code_ram_s1_address                           : out std_logic_vector(15 downto 0);                    -- address
			code_ram_s1_write                             : out std_logic;                                        -- write
			code_ram_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			code_ram_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			code_ram_s1_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			code_ram_s1_chipselect                        : out std_logic;                                        -- chipselect
			code_ram_s1_clken                             : out std_logic;                                        -- clken
			disp_7_seg_pio_disp_0_s1_address              : out std_logic_vector(1 downto 0);                     -- address
			disp_7_seg_pio_disp_0_s1_write                : out std_logic;                                        -- write
			disp_7_seg_pio_disp_0_s1_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			disp_7_seg_pio_disp_0_s1_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			disp_7_seg_pio_disp_0_s1_chipselect           : out std_logic;                                        -- chipselect
			disp_7_seg_pio_disp_1_s1_address              : out std_logic_vector(1 downto 0);                     -- address
			disp_7_seg_pio_disp_1_s1_write                : out std_logic;                                        -- write
			disp_7_seg_pio_disp_1_s1_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			disp_7_seg_pio_disp_1_s1_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			disp_7_seg_pio_disp_1_s1_chipselect           : out std_logic;                                        -- chipselect
			disp_7_seg_pio_disp_2_s1_address              : out std_logic_vector(1 downto 0);                     -- address
			disp_7_seg_pio_disp_2_s1_write                : out std_logic;                                        -- write
			disp_7_seg_pio_disp_2_s1_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			disp_7_seg_pio_disp_2_s1_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			disp_7_seg_pio_disp_2_s1_chipselect           : out std_logic;                                        -- chipselect
			disp_7_seg_pio_disp_3_s1_address              : out std_logic_vector(1 downto 0);                     -- address
			disp_7_seg_pio_disp_3_s1_write                : out std_logic;                                        -- write
			disp_7_seg_pio_disp_3_s1_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			disp_7_seg_pio_disp_3_s1_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			disp_7_seg_pio_disp_3_s1_chipselect           : out std_logic;                                        -- chipselect
			disp_7_seg_pio_disp_4_s1_address              : out std_logic_vector(1 downto 0);                     -- address
			disp_7_seg_pio_disp_4_s1_write                : out std_logic;                                        -- write
			disp_7_seg_pio_disp_4_s1_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			disp_7_seg_pio_disp_4_s1_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			disp_7_seg_pio_disp_4_s1_chipselect           : out std_logic;                                        -- chipselect
			disp_7_seg_pio_disp_5_s1_address              : out std_logic_vector(1 downto 0);                     -- address
			disp_7_seg_pio_disp_5_s1_write                : out std_logic;                                        -- write
			disp_7_seg_pio_disp_5_s1_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			disp_7_seg_pio_disp_5_s1_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			disp_7_seg_pio_disp_5_s1_chipselect           : out std_logic;                                        -- chipselect
			pio_leds_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			pio_leds_s1_write                             : out std_logic;                                        -- write
			pio_leds_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_leds_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_leds_s1_chipselect                        : out std_logic;                                        -- chipselect
			sdram_s1_address                              : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                : out std_logic;                                        -- write
			sdram_s1_read                                 : out std_logic;                                        -- read
			sdram_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                           : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                        : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                           : out std_logic;                                        -- chipselect
			timer_0_s1_address                            : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                              : out std_logic;                                        -- write
			timer_0_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                         : out std_logic                                         -- chipselect
		);
	end component system_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal altpll_0_c0_clk                                            : std_logic;                     -- altpll_0:c0 -> [sys_clk, av_dac:clk, av_uart:clk, av_vga:clk, code_ram:clk, disp_7_seg:pio_disp_0_clk_clk, disp_7_seg:pio_disp_1_clk_clk, disp_7_seg:pio_disp_2_clk_clk, disp_7_seg:pio_disp_3_clk_clk, disp_7_seg:pio_disp_4_clk_clk, disp_7_seg:pio_disp_5_clk_clk, mm_interconnect_0:altpll_0_c0_clk, pio_leds:clk, riscv_mk1_0:i_clk, rst_controller:clk, sdram:clk, timer_0:clk]
	signal riscv_mk1_0_avalon_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:riscv_mk1_0_avalon_master_waitrequest -> riscv_mk1_0:i_av_waitrequest
	signal riscv_mk1_0_avalon_master_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:riscv_mk1_0_avalon_master_readdata -> riscv_mk1_0:i_av_readdata
	signal riscv_mk1_0_avalon_master_address                          : std_logic_vector(29 downto 0); -- riscv_mk1_0:o_av_addr -> mm_interconnect_0:riscv_mk1_0_avalon_master_address
	signal riscv_mk1_0_avalon_master_byteenable                       : std_logic_vector(3 downto 0);  -- riscv_mk1_0:o_av_byteenable -> mm_interconnect_0:riscv_mk1_0_avalon_master_byteenable
	signal riscv_mk1_0_avalon_master_read                             : std_logic;                     -- riscv_mk1_0:o_av_read -> mm_interconnect_0:riscv_mk1_0_avalon_master_read
	signal riscv_mk1_0_avalon_master_write                            : std_logic;                     -- riscv_mk1_0:o_av_write -> mm_interconnect_0:riscv_mk1_0_avalon_master_write
	signal riscv_mk1_0_avalon_master_writedata                        : std_logic_vector(31 downto 0); -- riscv_mk1_0:o_av_writedata -> mm_interconnect_0:riscv_mk1_0_avalon_master_writedata
	signal mm_interconnect_0_av_dac_avalon_slave_chipselect           : std_logic;                     -- mm_interconnect_0:av_dac_avalon_slave_chipselect -> av_dac:avalon_chipselect
	signal mm_interconnect_0_av_dac_avalon_slave_readdata             : std_logic_vector(31 downto 0); -- av_dac:avalon_readdata -> mm_interconnect_0:av_dac_avalon_slave_readdata
	signal mm_interconnect_0_av_dac_avalon_slave_waitrequest          : std_logic;                     -- av_dac:avalon_waitrequest -> mm_interconnect_0:av_dac_avalon_slave_waitrequest
	signal mm_interconnect_0_av_dac_avalon_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:av_dac_avalon_slave_address -> av_dac:avalon_address
	signal mm_interconnect_0_av_dac_avalon_slave_read                 : std_logic;                     -- mm_interconnect_0:av_dac_avalon_slave_read -> av_dac:avalon_read
	signal mm_interconnect_0_av_dac_avalon_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:av_dac_avalon_slave_byteenable -> av_dac:avalon_byteenable
	signal mm_interconnect_0_av_dac_avalon_slave_write                : std_logic;                     -- mm_interconnect_0:av_dac_avalon_slave_write -> av_dac:avalon_write
	signal mm_interconnect_0_av_dac_avalon_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:av_dac_avalon_slave_writedata -> av_dac:avalon_writedata
	signal mm_interconnect_0_av_uart_avalon_slave_chipselect          : std_logic;                     -- mm_interconnect_0:av_uart_avalon_slave_chipselect -> av_uart:avalon_chipselect
	signal mm_interconnect_0_av_uart_avalon_slave_readdata            : std_logic_vector(31 downto 0); -- av_uart:avalon_readdata -> mm_interconnect_0:av_uart_avalon_slave_readdata
	signal mm_interconnect_0_av_uart_avalon_slave_waitrequest         : std_logic;                     -- av_uart:avalon_waitrequest -> mm_interconnect_0:av_uart_avalon_slave_waitrequest
	signal mm_interconnect_0_av_uart_avalon_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:av_uart_avalon_slave_address -> av_uart:avalon_address
	signal mm_interconnect_0_av_uart_avalon_slave_read                : std_logic;                     -- mm_interconnect_0:av_uart_avalon_slave_read -> av_uart:avalon_read
	signal mm_interconnect_0_av_uart_avalon_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:av_uart_avalon_slave_byteenable -> av_uart:avalon_byteenable
	signal mm_interconnect_0_av_uart_avalon_slave_write               : std_logic;                     -- mm_interconnect_0:av_uart_avalon_slave_write -> av_uart:avalon_write
	signal mm_interconnect_0_av_uart_avalon_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:av_uart_avalon_slave_writedata -> av_uart:avalon_writedata
	signal mm_interconnect_0_av_vga_avalon_slave_chipselect           : std_logic;                     -- mm_interconnect_0:av_vga_avalon_slave_chipselect -> av_vga:avalon_chipselect
	signal mm_interconnect_0_av_vga_avalon_slave_readdata             : std_logic_vector(31 downto 0); -- av_vga:avalon_readdata -> mm_interconnect_0:av_vga_avalon_slave_readdata
	signal mm_interconnect_0_av_vga_avalon_slave_waitrequest          : std_logic;                     -- av_vga:avalon_waitrequest -> mm_interconnect_0:av_vga_avalon_slave_waitrequest
	signal mm_interconnect_0_av_vga_avalon_slave_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:av_vga_avalon_slave_address -> av_vga:avalon_address
	signal mm_interconnect_0_av_vga_avalon_slave_read                 : std_logic;                     -- mm_interconnect_0:av_vga_avalon_slave_read -> av_vga:avalon_read
	signal mm_interconnect_0_av_vga_avalon_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:av_vga_avalon_slave_byteenable -> av_vga:avalon_byteenable
	signal mm_interconnect_0_av_vga_avalon_slave_write                : std_logic;                     -- mm_interconnect_0:av_vga_avalon_slave_write -> av_vga:avalon_write
	signal mm_interconnect_0_av_vga_avalon_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:av_vga_avalon_slave_writedata -> av_vga:avalon_writedata
	signal mm_interconnect_0_disp_7_seg_pio_disp_0_s1_chipselect      : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_0_s1_chipselect -> disp_7_seg:pio_disp_0_s1_chipselect
	signal mm_interconnect_0_disp_7_seg_pio_disp_0_s1_readdata        : std_logic_vector(31 downto 0); -- disp_7_seg:pio_disp_0_s1_readdata -> mm_interconnect_0:disp_7_seg_pio_disp_0_s1_readdata
	signal mm_interconnect_0_disp_7_seg_pio_disp_0_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:disp_7_seg_pio_disp_0_s1_address -> disp_7_seg:pio_disp_0_s1_address
	signal mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write           : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_0_s1_write -> mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write:in
	signal mm_interconnect_0_disp_7_seg_pio_disp_0_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:disp_7_seg_pio_disp_0_s1_writedata -> disp_7_seg:pio_disp_0_s1_writedata
	signal mm_interconnect_0_disp_7_seg_pio_disp_1_s1_chipselect      : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_1_s1_chipselect -> disp_7_seg:pio_disp_1_s1_chipselect
	signal mm_interconnect_0_disp_7_seg_pio_disp_1_s1_readdata        : std_logic_vector(31 downto 0); -- disp_7_seg:pio_disp_1_s1_readdata -> mm_interconnect_0:disp_7_seg_pio_disp_1_s1_readdata
	signal mm_interconnect_0_disp_7_seg_pio_disp_1_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:disp_7_seg_pio_disp_1_s1_address -> disp_7_seg:pio_disp_1_s1_address
	signal mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write           : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_1_s1_write -> mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write:in
	signal mm_interconnect_0_disp_7_seg_pio_disp_1_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:disp_7_seg_pio_disp_1_s1_writedata -> disp_7_seg:pio_disp_1_s1_writedata
	signal mm_interconnect_0_disp_7_seg_pio_disp_2_s1_chipselect      : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_2_s1_chipselect -> disp_7_seg:pio_disp_2_s1_chipselect
	signal mm_interconnect_0_disp_7_seg_pio_disp_2_s1_readdata        : std_logic_vector(31 downto 0); -- disp_7_seg:pio_disp_2_s1_readdata -> mm_interconnect_0:disp_7_seg_pio_disp_2_s1_readdata
	signal mm_interconnect_0_disp_7_seg_pio_disp_2_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:disp_7_seg_pio_disp_2_s1_address -> disp_7_seg:pio_disp_2_s1_address
	signal mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write           : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_2_s1_write -> mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write:in
	signal mm_interconnect_0_disp_7_seg_pio_disp_2_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:disp_7_seg_pio_disp_2_s1_writedata -> disp_7_seg:pio_disp_2_s1_writedata
	signal mm_interconnect_0_disp_7_seg_pio_disp_3_s1_chipselect      : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_3_s1_chipselect -> disp_7_seg:pio_disp_3_s1_chipselect
	signal mm_interconnect_0_disp_7_seg_pio_disp_3_s1_readdata        : std_logic_vector(31 downto 0); -- disp_7_seg:pio_disp_3_s1_readdata -> mm_interconnect_0:disp_7_seg_pio_disp_3_s1_readdata
	signal mm_interconnect_0_disp_7_seg_pio_disp_3_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:disp_7_seg_pio_disp_3_s1_address -> disp_7_seg:pio_disp_3_s1_address
	signal mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write           : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_3_s1_write -> mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write:in
	signal mm_interconnect_0_disp_7_seg_pio_disp_3_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:disp_7_seg_pio_disp_3_s1_writedata -> disp_7_seg:pio_disp_3_s1_writedata
	signal mm_interconnect_0_disp_7_seg_pio_disp_4_s1_chipselect      : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_4_s1_chipselect -> disp_7_seg:pio_disp_4_s1_chipselect
	signal mm_interconnect_0_disp_7_seg_pio_disp_4_s1_readdata        : std_logic_vector(31 downto 0); -- disp_7_seg:pio_disp_4_s1_readdata -> mm_interconnect_0:disp_7_seg_pio_disp_4_s1_readdata
	signal mm_interconnect_0_disp_7_seg_pio_disp_4_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:disp_7_seg_pio_disp_4_s1_address -> disp_7_seg:pio_disp_4_s1_address
	signal mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write           : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_4_s1_write -> mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write:in
	signal mm_interconnect_0_disp_7_seg_pio_disp_4_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:disp_7_seg_pio_disp_4_s1_writedata -> disp_7_seg:pio_disp_4_s1_writedata
	signal mm_interconnect_0_disp_7_seg_pio_disp_5_s1_chipselect      : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_5_s1_chipselect -> disp_7_seg:pio_disp_5_s1_chipselect
	signal mm_interconnect_0_disp_7_seg_pio_disp_5_s1_readdata        : std_logic_vector(31 downto 0); -- disp_7_seg:pio_disp_5_s1_readdata -> mm_interconnect_0:disp_7_seg_pio_disp_5_s1_readdata
	signal mm_interconnect_0_disp_7_seg_pio_disp_5_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:disp_7_seg_pio_disp_5_s1_address -> disp_7_seg:pio_disp_5_s1_address
	signal mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write           : std_logic;                     -- mm_interconnect_0:disp_7_seg_pio_disp_5_s1_write -> mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write:in
	signal mm_interconnect_0_disp_7_seg_pio_disp_5_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:disp_7_seg_pio_disp_5_s1_writedata -> disp_7_seg:pio_disp_5_s1_writedata
	signal mm_interconnect_0_code_ram_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:code_ram_s1_chipselect -> code_ram:chipselect
	signal mm_interconnect_0_code_ram_s1_readdata                     : std_logic_vector(31 downto 0); -- code_ram:readdata -> mm_interconnect_0:code_ram_s1_readdata
	signal mm_interconnect_0_code_ram_s1_address                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:code_ram_s1_address -> code_ram:address
	signal mm_interconnect_0_code_ram_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:code_ram_s1_byteenable -> code_ram:byteenable
	signal mm_interconnect_0_code_ram_s1_write                        : std_logic;                     -- mm_interconnect_0:code_ram_s1_write -> code_ram:write
	signal mm_interconnect_0_code_ram_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:code_ram_s1_writedata -> code_ram:writedata
	signal mm_interconnect_0_code_ram_s1_clken                        : std_logic;                     -- mm_interconnect_0:code_ram_s1_clken -> code_ram:clken
	signal mm_interconnect_0_pio_leds_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:pio_leds_s1_chipselect -> pio_leds:chipselect
	signal mm_interconnect_0_pio_leds_s1_readdata                     : std_logic_vector(31 downto 0); -- pio_leds:readdata -> mm_interconnect_0:pio_leds_s1_readdata
	signal mm_interconnect_0_pio_leds_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_leds_s1_address -> pio_leds:address
	signal mm_interconnect_0_pio_leds_s1_write                        : std_logic;                     -- mm_interconnect_0:pio_leds_s1_write -> mm_interconnect_0_pio_leds_s1_write:in
	signal mm_interconnect_0_pio_leds_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_leds_s1_writedata -> pio_leds:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                        : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                     : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                         : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                            : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                   : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                           : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_timer_0_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                      : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                         : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal rst_controller_reset_out_reset                             : std_logic;                     -- rst_controller:reset_out -> [av_dac:reset, av_uart:reset, av_vga:reset, code_ram:reset, mm_interconnect_0:riscv_mk1_0_reset_reset_bridge_in_reset_reset, riscv_mk1_0:i_rst, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                         : std_logic;                     -- rst_controller:reset_req -> [code_ram:reset_req, rst_translator:reset_req_in]
	signal rst_reset_n_ports_inv                                      : std_logic;                     -- rst_reset_n:inv -> [altpll_0:reset, rst_controller:reset_in0]
	signal mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write:inv -> disp_7_seg:pio_disp_0_s1_write_n
	signal mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write:inv -> disp_7_seg:pio_disp_1_s1_write_n
	signal mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write:inv -> disp_7_seg:pio_disp_2_s1_write_n
	signal mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write:inv -> disp_7_seg:pio_disp_3_s1_write_n
	signal mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write:inv -> disp_7_seg:pio_disp_4_s1_write_n
	signal mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write:inv -> disp_7_seg:pio_disp_5_s1_write_n
	signal mm_interconnect_0_pio_leds_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_pio_leds_s1_write:inv -> pio_leds:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                  : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv            : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_reset_out_reset:inv -> [disp_7_seg:pio_disp_0_reset_reset_n, disp_7_seg:pio_disp_1_reset_reset_n, disp_7_seg:pio_disp_2_reset_reset_n, disp_7_seg:pio_disp_3_reset_reset_n, disp_7_seg:pio_disp_4_reset_reset_n, disp_7_seg:pio_disp_5_reset_reset_n, pio_leds:reset_n, sdram:reset_n, timer_0:reset_n]

begin

	altpll_0 : component system_altpll_0
		port map (
			clk                => clk_clk,               --       inclk_interface.clk
			reset              => rst_reset_n_ports_inv, -- inclk_interface_reset.reset
			read               => open,                  --             pll_slave.read
			write              => open,                  --                      .write
			address            => open,                  --                      .address
			readdata           => open,                  --                      .readdata
			writedata          => open,                  --                      .writedata
			c0                 => altpll_0_c0_clk,       --                    c0.clk
			c1                 => clk_sdram_clk,         --                    c1.clk
			scandone           => open,                  --           (terminated)
			scandataout        => open,                  --           (terminated)
			c2                 => open,                  --           (terminated)
			c3                 => open,                  --           (terminated)
			c4                 => open,                  --           (terminated)
			areset             => '0',                   --           (terminated)
			locked             => open,                  --           (terminated)
			phasedone          => open,                  --           (terminated)
			phasecounterselect => "000",                 --           (terminated)
			phaseupdown        => '0',                   --           (terminated)
			phasestep          => '0',                   --           (terminated)
			scanclk            => '0',                   --           (terminated)
			scanclkena         => '0',                   --           (terminated)
			scandata           => '0',                   --           (terminated)
			configupdate       => '0'                    --           (terminated)
		);

	av_dac : component system_av_dac
		port map (
			clk                => altpll_0_c0_clk,                                   --                clk.clk
			reset              => rst_controller_reset_out_reset,                    --              reset.reset
			avalon_address     => mm_interconnect_0_av_dac_avalon_slave_address(0),  --       avalon_slave.address
			avalon_byteenable  => mm_interconnect_0_av_dac_avalon_slave_byteenable,  --                   .byteenable
			avalon_chipselect  => mm_interconnect_0_av_dac_avalon_slave_chipselect,  --                   .chipselect
			avalon_read        => mm_interconnect_0_av_dac_avalon_slave_read,        --                   .read
			avalon_write       => mm_interconnect_0_av_dac_avalon_slave_write,       --                   .write
			avalon_writedata   => mm_interconnect_0_av_dac_avalon_slave_writedata,   --                   .writedata
			avalon_readdata    => mm_interconnect_0_av_dac_avalon_slave_readdata,    --                   .readdata
			avalon_waitrequest => mm_interconnect_0_av_dac_avalon_slave_waitrequest, --                   .waitrequest
			avalon_irq         => open,                                              --          interrupt.irq
			acknowledge        => av_dac_external_interface_acknowledge,             -- external_interface.export
			irq                => av_dac_external_interface_irq,                     --                   .export
			address            => av_dac_external_interface_address,                 --                   .export
			bus_enable         => av_dac_external_interface_bus_enable,              --                   .export
			byte_enable        => av_dac_external_interface_byte_enable,             --                   .export
			rw                 => av_dac_external_interface_rw,                      --                   .export
			write_data         => av_dac_external_interface_write_data,              --                   .export
			read_data          => av_dac_external_interface_read_data                --                   .export
		);

	av_uart : component system_av_dac
		port map (
			clk                => altpll_0_c0_clk,                                    --                clk.clk
			reset              => rst_controller_reset_out_reset,                     --              reset.reset
			avalon_address     => mm_interconnect_0_av_uart_avalon_slave_address(0),  --       avalon_slave.address
			avalon_byteenable  => mm_interconnect_0_av_uart_avalon_slave_byteenable,  --                   .byteenable
			avalon_chipselect  => mm_interconnect_0_av_uart_avalon_slave_chipselect,  --                   .chipselect
			avalon_read        => mm_interconnect_0_av_uart_avalon_slave_read,        --                   .read
			avalon_write       => mm_interconnect_0_av_uart_avalon_slave_write,       --                   .write
			avalon_writedata   => mm_interconnect_0_av_uart_avalon_slave_writedata,   --                   .writedata
			avalon_readdata    => mm_interconnect_0_av_uart_avalon_slave_readdata,    --                   .readdata
			avalon_waitrequest => mm_interconnect_0_av_uart_avalon_slave_waitrequest, --                   .waitrequest
			avalon_irq         => open,                                               --          interrupt.irq
			acknowledge        => av_uart_external_interface_acknowledge,             -- external_interface.export
			irq                => av_uart_external_interface_irq,                     --                   .export
			address            => av_uart_external_interface_address,                 --                   .export
			bus_enable         => av_uart_external_interface_bus_enable,              --                   .export
			byte_enable        => av_uart_external_interface_byte_enable,             --                   .export
			rw                 => av_uart_external_interface_rw,                      --                   .export
			write_data         => av_uart_external_interface_write_data,              --                   .export
			read_data          => av_uart_external_interface_read_data                --                   .export
		);

	av_vga : component system_av_vga
		port map (
			clk                => altpll_0_c0_clk,                                   --                clk.clk
			reset              => rst_controller_reset_out_reset,                    --              reset.reset
			avalon_address     => mm_interconnect_0_av_vga_avalon_slave_address,     --       avalon_slave.address
			avalon_byteenable  => mm_interconnect_0_av_vga_avalon_slave_byteenable,  --                   .byteenable
			avalon_chipselect  => mm_interconnect_0_av_vga_avalon_slave_chipselect,  --                   .chipselect
			avalon_read        => mm_interconnect_0_av_vga_avalon_slave_read,        --                   .read
			avalon_write       => mm_interconnect_0_av_vga_avalon_slave_write,       --                   .write
			avalon_writedata   => mm_interconnect_0_av_vga_avalon_slave_writedata,   --                   .writedata
			avalon_readdata    => mm_interconnect_0_av_vga_avalon_slave_readdata,    --                   .readdata
			avalon_waitrequest => mm_interconnect_0_av_vga_avalon_slave_waitrequest, --                   .waitrequest
			avalon_irq         => open,                                              --          interrupt.irq
			acknowledge        => av_vga_external_interface_acknowledge,             -- external_interface.export
			irq                => av_vga_external_interface_irq,                     --                   .export
			address            => av_vga_external_interface_address,                 --                   .export
			bus_enable         => av_vga_external_interface_bus_enable,              --                   .export
			byte_enable        => av_vga_external_interface_byte_enable,             --                   .export
			rw                 => av_vga_external_interface_rw,                      --                   .export
			write_data         => av_vga_external_interface_write_data,              --                   .export
			read_data          => av_vga_external_interface_read_data                --                   .export
		);

	code_ram : component system_code_ram
		port map (
			clk        => altpll_0_c0_clk,                          --   clk1.clk
			address    => mm_interconnect_0_code_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_code_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_code_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_code_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_code_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_code_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_code_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,           -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,       --       .reset_req
			freeze     => '0'                                       -- (terminated)
		);

	disp_7_seg : component system_disp_7_seg
		port map (
			pio_disp_0_clk_clk                    => altpll_0_c0_clk,                                            --                 pio_disp_0_clk.clk
			pio_disp_0_external_connection_export => disp0_export,                                               -- pio_disp_0_external_connection.export
			pio_disp_0_reset_reset_n              => rst_controller_reset_out_reset_ports_inv,                   --               pio_disp_0_reset.reset_n
			pio_disp_0_s1_address                 => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_address,         --                  pio_disp_0_s1.address
			pio_disp_0_s1_write_n                 => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write_ports_inv, --                               .write_n
			pio_disp_0_s1_writedata               => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_writedata,       --                               .writedata
			pio_disp_0_s1_chipselect              => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_chipselect,      --                               .chipselect
			pio_disp_0_s1_readdata                => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_readdata,        --                               .readdata
			pio_disp_1_clk_clk                    => altpll_0_c0_clk,                                            --                 pio_disp_1_clk.clk
			pio_disp_1_external_connection_export => disp1_export,                                               -- pio_disp_1_external_connection.export
			pio_disp_1_reset_reset_n              => rst_controller_reset_out_reset_ports_inv,                   --               pio_disp_1_reset.reset_n
			pio_disp_1_s1_address                 => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_address,         --                  pio_disp_1_s1.address
			pio_disp_1_s1_write_n                 => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write_ports_inv, --                               .write_n
			pio_disp_1_s1_writedata               => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_writedata,       --                               .writedata
			pio_disp_1_s1_chipselect              => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_chipselect,      --                               .chipselect
			pio_disp_1_s1_readdata                => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_readdata,        --                               .readdata
			pio_disp_2_clk_clk                    => altpll_0_c0_clk,                                            --                 pio_disp_2_clk.clk
			pio_disp_2_external_connection_export => disp2_export,                                               -- pio_disp_2_external_connection.export
			pio_disp_2_reset_reset_n              => rst_controller_reset_out_reset_ports_inv,                   --               pio_disp_2_reset.reset_n
			pio_disp_2_s1_address                 => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_address,         --                  pio_disp_2_s1.address
			pio_disp_2_s1_write_n                 => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write_ports_inv, --                               .write_n
			pio_disp_2_s1_writedata               => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_writedata,       --                               .writedata
			pio_disp_2_s1_chipselect              => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_chipselect,      --                               .chipselect
			pio_disp_2_s1_readdata                => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_readdata,        --                               .readdata
			pio_disp_3_clk_clk                    => altpll_0_c0_clk,                                            --                 pio_disp_3_clk.clk
			pio_disp_3_external_connection_export => disp3_export,                                               -- pio_disp_3_external_connection.export
			pio_disp_3_reset_reset_n              => rst_controller_reset_out_reset_ports_inv,                   --               pio_disp_3_reset.reset_n
			pio_disp_3_s1_address                 => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_address,         --                  pio_disp_3_s1.address
			pio_disp_3_s1_write_n                 => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write_ports_inv, --                               .write_n
			pio_disp_3_s1_writedata               => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_writedata,       --                               .writedata
			pio_disp_3_s1_chipselect              => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_chipselect,      --                               .chipselect
			pio_disp_3_s1_readdata                => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_readdata,        --                               .readdata
			pio_disp_4_clk_clk                    => altpll_0_c0_clk,                                            --                 pio_disp_4_clk.clk
			pio_disp_4_external_connection_export => disp4_export,                                               -- pio_disp_4_external_connection.export
			pio_disp_4_reset_reset_n              => rst_controller_reset_out_reset_ports_inv,                   --               pio_disp_4_reset.reset_n
			pio_disp_4_s1_address                 => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_address,         --                  pio_disp_4_s1.address
			pio_disp_4_s1_write_n                 => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write_ports_inv, --                               .write_n
			pio_disp_4_s1_writedata               => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_writedata,       --                               .writedata
			pio_disp_4_s1_chipselect              => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_chipselect,      --                               .chipselect
			pio_disp_4_s1_readdata                => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_readdata,        --                               .readdata
			pio_disp_5_clk_clk                    => altpll_0_c0_clk,                                            --                 pio_disp_5_clk.clk
			pio_disp_5_external_connection_export => disp5_export,                                               -- pio_disp_5_external_connection.export
			pio_disp_5_reset_reset_n              => rst_controller_reset_out_reset_ports_inv,                   --               pio_disp_5_reset.reset_n
			pio_disp_5_s1_address                 => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_address,         --                  pio_disp_5_s1.address
			pio_disp_5_s1_write_n                 => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write_ports_inv, --                               .write_n
			pio_disp_5_s1_writedata               => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_writedata,       --                               .writedata
			pio_disp_5_s1_chipselect              => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_chipselect,      --                               .chipselect
			pio_disp_5_s1_readdata                => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_readdata         --                               .readdata
		);

	pio_leds : component system_pio_leds
		port map (
			clk        => altpll_0_c0_clk,                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_leds_s1_readdata,        --                    .readdata
			out_port   => leds_export                                    -- external_connection.export
		);

	riscv_mk1_0 : component riscv_mk1
		port map (
			o_av_addr        => riscv_mk1_0_avalon_master_address,     -- avalon_master.address
			o_av_byteenable  => riscv_mk1_0_avalon_master_byteenable,  --              .byteenable
			o_av_read        => riscv_mk1_0_avalon_master_read,        --              .read
			o_av_write       => riscv_mk1_0_avalon_master_write,       --              .write
			i_av_waitrequest => riscv_mk1_0_avalon_master_waitrequest, --              .waitrequest
			o_av_writedata   => riscv_mk1_0_avalon_master_writedata,   --              .writedata
			i_av_readdata    => riscv_mk1_0_avalon_master_readdata,    --              .readdata
			i_clk            => altpll_0_c0_clk,                       --         clock.clk
			i_rst            => rst_controller_reset_out_reset         --         reset.reset
		);

	sdram : component system_sdram
		port map (
			clk            => altpll_0_c0_clk,                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	timer_0 : component system_timer_0
		port map (
			clk        => altpll_0_c0_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => open                                          --   irq.irq
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			altpll_0_c0_clk                               => altpll_0_c0_clk,                                       --                             altpll_0_c0.clk
			riscv_mk1_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                        -- riscv_mk1_0_reset_reset_bridge_in_reset.reset
			riscv_mk1_0_avalon_master_address             => riscv_mk1_0_avalon_master_address,                     --               riscv_mk1_0_avalon_master.address
			riscv_mk1_0_avalon_master_waitrequest         => riscv_mk1_0_avalon_master_waitrequest,                 --                                        .waitrequest
			riscv_mk1_0_avalon_master_byteenable          => riscv_mk1_0_avalon_master_byteenable,                  --                                        .byteenable
			riscv_mk1_0_avalon_master_read                => riscv_mk1_0_avalon_master_read,                        --                                        .read
			riscv_mk1_0_avalon_master_readdata            => riscv_mk1_0_avalon_master_readdata,                    --                                        .readdata
			riscv_mk1_0_avalon_master_write               => riscv_mk1_0_avalon_master_write,                       --                                        .write
			riscv_mk1_0_avalon_master_writedata           => riscv_mk1_0_avalon_master_writedata,                   --                                        .writedata
			av_dac_avalon_slave_address                   => mm_interconnect_0_av_dac_avalon_slave_address,         --                     av_dac_avalon_slave.address
			av_dac_avalon_slave_write                     => mm_interconnect_0_av_dac_avalon_slave_write,           --                                        .write
			av_dac_avalon_slave_read                      => mm_interconnect_0_av_dac_avalon_slave_read,            --                                        .read
			av_dac_avalon_slave_readdata                  => mm_interconnect_0_av_dac_avalon_slave_readdata,        --                                        .readdata
			av_dac_avalon_slave_writedata                 => mm_interconnect_0_av_dac_avalon_slave_writedata,       --                                        .writedata
			av_dac_avalon_slave_byteenable                => mm_interconnect_0_av_dac_avalon_slave_byteenable,      --                                        .byteenable
			av_dac_avalon_slave_waitrequest               => mm_interconnect_0_av_dac_avalon_slave_waitrequest,     --                                        .waitrequest
			av_dac_avalon_slave_chipselect                => mm_interconnect_0_av_dac_avalon_slave_chipselect,      --                                        .chipselect
			av_uart_avalon_slave_address                  => mm_interconnect_0_av_uart_avalon_slave_address,        --                    av_uart_avalon_slave.address
			av_uart_avalon_slave_write                    => mm_interconnect_0_av_uart_avalon_slave_write,          --                                        .write
			av_uart_avalon_slave_read                     => mm_interconnect_0_av_uart_avalon_slave_read,           --                                        .read
			av_uart_avalon_slave_readdata                 => mm_interconnect_0_av_uart_avalon_slave_readdata,       --                                        .readdata
			av_uart_avalon_slave_writedata                => mm_interconnect_0_av_uart_avalon_slave_writedata,      --                                        .writedata
			av_uart_avalon_slave_byteenable               => mm_interconnect_0_av_uart_avalon_slave_byteenable,     --                                        .byteenable
			av_uart_avalon_slave_waitrequest              => mm_interconnect_0_av_uart_avalon_slave_waitrequest,    --                                        .waitrequest
			av_uart_avalon_slave_chipselect               => mm_interconnect_0_av_uart_avalon_slave_chipselect,     --                                        .chipselect
			av_vga_avalon_slave_address                   => mm_interconnect_0_av_vga_avalon_slave_address,         --                     av_vga_avalon_slave.address
			av_vga_avalon_slave_write                     => mm_interconnect_0_av_vga_avalon_slave_write,           --                                        .write
			av_vga_avalon_slave_read                      => mm_interconnect_0_av_vga_avalon_slave_read,            --                                        .read
			av_vga_avalon_slave_readdata                  => mm_interconnect_0_av_vga_avalon_slave_readdata,        --                                        .readdata
			av_vga_avalon_slave_writedata                 => mm_interconnect_0_av_vga_avalon_slave_writedata,       --                                        .writedata
			av_vga_avalon_slave_byteenable                => mm_interconnect_0_av_vga_avalon_slave_byteenable,      --                                        .byteenable
			av_vga_avalon_slave_waitrequest               => mm_interconnect_0_av_vga_avalon_slave_waitrequest,     --                                        .waitrequest
			av_vga_avalon_slave_chipselect                => mm_interconnect_0_av_vga_avalon_slave_chipselect,      --                                        .chipselect
			code_ram_s1_address                           => mm_interconnect_0_code_ram_s1_address,                 --                             code_ram_s1.address
			code_ram_s1_write                             => mm_interconnect_0_code_ram_s1_write,                   --                                        .write
			code_ram_s1_readdata                          => mm_interconnect_0_code_ram_s1_readdata,                --                                        .readdata
			code_ram_s1_writedata                         => mm_interconnect_0_code_ram_s1_writedata,               --                                        .writedata
			code_ram_s1_byteenable                        => mm_interconnect_0_code_ram_s1_byteenable,              --                                        .byteenable
			code_ram_s1_chipselect                        => mm_interconnect_0_code_ram_s1_chipselect,              --                                        .chipselect
			code_ram_s1_clken                             => mm_interconnect_0_code_ram_s1_clken,                   --                                        .clken
			disp_7_seg_pio_disp_0_s1_address              => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_address,    --                disp_7_seg_pio_disp_0_s1.address
			disp_7_seg_pio_disp_0_s1_write                => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write,      --                                        .write
			disp_7_seg_pio_disp_0_s1_readdata             => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_readdata,   --                                        .readdata
			disp_7_seg_pio_disp_0_s1_writedata            => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_writedata,  --                                        .writedata
			disp_7_seg_pio_disp_0_s1_chipselect           => mm_interconnect_0_disp_7_seg_pio_disp_0_s1_chipselect, --                                        .chipselect
			disp_7_seg_pio_disp_1_s1_address              => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_address,    --                disp_7_seg_pio_disp_1_s1.address
			disp_7_seg_pio_disp_1_s1_write                => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write,      --                                        .write
			disp_7_seg_pio_disp_1_s1_readdata             => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_readdata,   --                                        .readdata
			disp_7_seg_pio_disp_1_s1_writedata            => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_writedata,  --                                        .writedata
			disp_7_seg_pio_disp_1_s1_chipselect           => mm_interconnect_0_disp_7_seg_pio_disp_1_s1_chipselect, --                                        .chipselect
			disp_7_seg_pio_disp_2_s1_address              => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_address,    --                disp_7_seg_pio_disp_2_s1.address
			disp_7_seg_pio_disp_2_s1_write                => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write,      --                                        .write
			disp_7_seg_pio_disp_2_s1_readdata             => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_readdata,   --                                        .readdata
			disp_7_seg_pio_disp_2_s1_writedata            => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_writedata,  --                                        .writedata
			disp_7_seg_pio_disp_2_s1_chipselect           => mm_interconnect_0_disp_7_seg_pio_disp_2_s1_chipselect, --                                        .chipselect
			disp_7_seg_pio_disp_3_s1_address              => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_address,    --                disp_7_seg_pio_disp_3_s1.address
			disp_7_seg_pio_disp_3_s1_write                => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write,      --                                        .write
			disp_7_seg_pio_disp_3_s1_readdata             => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_readdata,   --                                        .readdata
			disp_7_seg_pio_disp_3_s1_writedata            => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_writedata,  --                                        .writedata
			disp_7_seg_pio_disp_3_s1_chipselect           => mm_interconnect_0_disp_7_seg_pio_disp_3_s1_chipselect, --                                        .chipselect
			disp_7_seg_pio_disp_4_s1_address              => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_address,    --                disp_7_seg_pio_disp_4_s1.address
			disp_7_seg_pio_disp_4_s1_write                => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write,      --                                        .write
			disp_7_seg_pio_disp_4_s1_readdata             => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_readdata,   --                                        .readdata
			disp_7_seg_pio_disp_4_s1_writedata            => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_writedata,  --                                        .writedata
			disp_7_seg_pio_disp_4_s1_chipselect           => mm_interconnect_0_disp_7_seg_pio_disp_4_s1_chipselect, --                                        .chipselect
			disp_7_seg_pio_disp_5_s1_address              => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_address,    --                disp_7_seg_pio_disp_5_s1.address
			disp_7_seg_pio_disp_5_s1_write                => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write,      --                                        .write
			disp_7_seg_pio_disp_5_s1_readdata             => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_readdata,   --                                        .readdata
			disp_7_seg_pio_disp_5_s1_writedata            => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_writedata,  --                                        .writedata
			disp_7_seg_pio_disp_5_s1_chipselect           => mm_interconnect_0_disp_7_seg_pio_disp_5_s1_chipselect, --                                        .chipselect
			pio_leds_s1_address                           => mm_interconnect_0_pio_leds_s1_address,                 --                             pio_leds_s1.address
			pio_leds_s1_write                             => mm_interconnect_0_pio_leds_s1_write,                   --                                        .write
			pio_leds_s1_readdata                          => mm_interconnect_0_pio_leds_s1_readdata,                --                                        .readdata
			pio_leds_s1_writedata                         => mm_interconnect_0_pio_leds_s1_writedata,               --                                        .writedata
			pio_leds_s1_chipselect                        => mm_interconnect_0_pio_leds_s1_chipselect,              --                                        .chipselect
			sdram_s1_address                              => mm_interconnect_0_sdram_s1_address,                    --                                sdram_s1.address
			sdram_s1_write                                => mm_interconnect_0_sdram_s1_write,                      --                                        .write
			sdram_s1_read                                 => mm_interconnect_0_sdram_s1_read,                       --                                        .read
			sdram_s1_readdata                             => mm_interconnect_0_sdram_s1_readdata,                   --                                        .readdata
			sdram_s1_writedata                            => mm_interconnect_0_sdram_s1_writedata,                  --                                        .writedata
			sdram_s1_byteenable                           => mm_interconnect_0_sdram_s1_byteenable,                 --                                        .byteenable
			sdram_s1_readdatavalid                        => mm_interconnect_0_sdram_s1_readdatavalid,              --                                        .readdatavalid
			sdram_s1_waitrequest                          => mm_interconnect_0_sdram_s1_waitrequest,                --                                        .waitrequest
			sdram_s1_chipselect                           => mm_interconnect_0_sdram_s1_chipselect,                 --                                        .chipselect
			timer_0_s1_address                            => mm_interconnect_0_timer_0_s1_address,                  --                              timer_0_s1.address
			timer_0_s1_write                              => mm_interconnect_0_timer_0_s1_write,                    --                                        .write
			timer_0_s1_readdata                           => mm_interconnect_0_timer_0_s1_readdata,                 --                                        .readdata
			timer_0_s1_writedata                          => mm_interconnect_0_timer_0_s1_writedata,                --                                        .writedata
			timer_0_s1_chipselect                         => mm_interconnect_0_timer_0_s1_chipselect                --                                        .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => altpll_0_c0_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_reset_n_ports_inv <= not rst_reset_n;

	mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write_ports_inv <= not mm_interconnect_0_disp_7_seg_pio_disp_0_s1_write;

	mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write_ports_inv <= not mm_interconnect_0_disp_7_seg_pio_disp_1_s1_write;

	mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write_ports_inv <= not mm_interconnect_0_disp_7_seg_pio_disp_2_s1_write;

	mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write_ports_inv <= not mm_interconnect_0_disp_7_seg_pio_disp_3_s1_write;

	mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write_ports_inv <= not mm_interconnect_0_disp_7_seg_pio_disp_4_s1_write;

	mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write_ports_inv <= not mm_interconnect_0_disp_7_seg_pio_disp_5_s1_write;

	mm_interconnect_0_pio_leds_s1_write_ports_inv <= not mm_interconnect_0_pio_leds_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	sys_clk <= altpll_0_c0_clk;

end architecture rtl; -- of system
