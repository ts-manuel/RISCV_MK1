00021197
2b018193
08000117
ff810113
00018297
25c28293
04000317
fe830313
04007397
66038393
406383b3
00038e63
0002ae03
01c32023
00428293
00430313
ffc38393
fe9ff06f
04007297
6ec28293
04007317
74430313
40530333
00030a63
0002a023
00428293
ffc30313
ff1ff06f
0040006f
00021197
23c18193
04007517
60450513
04007617
71060613
40a60633
00000593
36c040ef
00012517
be450513
00050863
00008517
be050513
3d1110ef
2c4040ef
00012503
00410593
00000613
739170ef
27c0406f
ff010113
00812423
04007437
73444783
00112623
02079263
00000793
00078a63
04007537
68050513
00000097
000000e7
00100793
72f40a23
00c12083
00812403
01010113
00008067
00000793
00078e63
040075b7
04007537
73858593
68050513
00000317
00000067
00008067
04007737
77872783
00078a63
00a78533
76a72c23
00078513
00008067
040077b7
79478793
00a78533
76a72c23
00078513
00008067
fd010113
01712623
02112623
02812423
02912223
03212023
01312e23
01412c23
01512a23
01612823
01812423
00b50bb3
09757863
00020a37
00050b13
01050913
00020c37
00020ab7
b1da0a13
000209b7
000b0593
78cc0513
000b0493
358040ef
000b0413
00044583
794a8513
00140413
344040ef
fe8918e3
02000513
390040ef
0004c703
79c98513
02e00593
00ea07b3
0007c783
0977f793
04078c63
00148493
00070593
310040ef
fc991ce3
00a00513
010b0b13
358040ef
01090913
f97b6ae3
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
00148493
79c98513
2bc040ef
f89912e3
00a00513
010b0b13
304040ef
01090913
f57b60e3
fadff06f
040077b7
77c7c703
00100513
02071063
20000737
00072703
040076b7
00f75513
00157513
76e68ea3
76a78e23
00008067
04007737
77c74783
00078a63
040077b7
77d7c503
76070e23
00008067
040075b7
20000637
000086b7
00062783
0ff7f513
76a58ea3
00d7f7b3
fe0788e3
fd9ff06f
20000737
04000693
00472783
0107d793
fed79ce3
00a70023
00008067
00060513
02c05663
00c588b3
20000737
04000693
0005c803
00158593
00472783
0107d793
fed79ce3
01070023
feb894e3
00008067
00060513
06c05463
04007637
77c64783
00a58333
040076b7
200008b7
00008837
0140006f
77d6c703
fee58fa3
00000793
02658c63
00158593
fe0796e3
0008a783
0ff7f713
76e68ea3
0107f7b3
fc079ee3
0008a783
0ff7f713
76e68ea3
0107f7b3
fc078ee3
fc5ff06f
76060e23
00008067
f8010113
05712e23
02050b93
06812c23
06112e23
06912a23
07212823
07312623
07412423
07512223
07612023
05812c23
05912a23
05a12823
05b12623
00050413
00a12823
01712623
00042503
000214b7
00440413
495030ef
a404a583
438030ef
00050c13
07c42503
481030ef
a404a583
424030ef
00050c93
03c42503
46d030ef
000217b7
a447a583
40c030ef
00050a93
0bc42503
455030ef
000217b7
a487a583
3f4030ef
00050b93
09c42503
43d030ef
000217b7
a4c7a583
3dc030ef
00050493
01c42503
425030ef
000217b7
a507a583
3c4030ef
00050a13
0dc42503
40d030ef
000217b7
a547a583
3ac030ef
00050d13
05c42503
3f5030ef
000217b7
a587a583
394030ef
00050993
00050593
00048513
6fc030ef
00050b13
000d0593
000a0513
721020ef
00050913
000d0593
000a0513
6dc030ef
00050d93
00098593
00048513
701020ef
00050a13
000b8593
000a8513
6f1020ef
00050993
000a0593
00090513
6e1020ef
00050493
000d8593
000b0513
6d1020ef
000217b7
a5c7a583
318030ef
00050d13
000c8593
000c0513
6b5020ef
00050693
000c8593
000c0513
00068c93
66c030ef
00050c13
000b8593
000a8513
65c030ef
00021bb7
a60ba583
2d8030ef
00098593
648030ef
000217b7
a647a583
00050a93
000d8513
2bc030ef
000d0593
62c030ef
00050d93
000a0593
00090513
61c030ef
a60ba583
29c030ef
00048593
641020ef
000d8593
604030ef
00050913
000c8593
00098513
629020ef
00050a13
000a8593
000c0513
619020ef
00050713
000a8593
000c0513
00070a93
5d0030ef
00050c13
00098593
000c8513
5c0030ef
000217b7
a687a583
00050c93
000b0513
234030ef
000d0593
5d9020ef
00090593
59c030ef
00050d13
00048593
000d8513
58c030ef
00050993
000a0593
00048513
5b1020ef
1e5030ef
00098593
fea42e23
000a8513
59d020ef
1d1030ef
000c0593
00a42e23
00090513
589020ef
1bd030ef
000d0593
02a42e23
000c8513
575020ef
1a9030ef
000d0593
04a42e23
000c8513
52c030ef
195030ef
00090593
06a42e23
000c0513
518030ef
181030ef
00098593
08a42e23
000a8513
504030ef
16d030ef
00048593
0aa42e23
000a0513
4f0030ef
159030ef
00c12783
0ca42e23
d0879ee3
00078b93
000217b7
a407a783
01012b03
000b8c93
00f12c23
000217b7
a447a783
00f12e23
000217b7
a487a783
02f12023
000217b7
a4c7a783
02f12223
000217b7
a507a783
02f12423
000217b7
a547a783
02f12623
000217b7
a587a783
02f12823
000217b7
a5c7a783
02f12a23
000217b7
a607a783
00f12623
000217b7
a647a783
02f12c23
000217b7
a687a783
02f12e23
100b0793
00f12a23
0080006f
020c8c93
000b2503
115030ef
01812403
00040593
0b4030ef
00050a93
010b2503
0fd030ef
00040593
0a0030ef
00050c13
008b2503
0e9030ef
01c12583
08c030ef
00050a13
018b2503
0d5030ef
02012583
078030ef
00050713
014b2503
00e12823
0bd030ef
02412583
060030ef
00050413
004b2503
0a9030ef
02812583
04c030ef
00050993
01cb2503
095030ef
02c12583
038030ef
00050d13
00cb2503
081030ef
03012583
024030ef
00050913
00050593
00040513
38c030ef
00050b93
000d0593
00098513
3b1020ef
00050493
000d0593
00098513
36c030ef
00050d93
00090593
00040513
391020ef
01012703
00050993
000a0513
00070593
37d020ef
00050913
00098593
00048513
36d020ef
00050413
000d8593
000b8513
35d020ef
03412583
7a9020ef
00050d13
000c0593
000a8513
345020ef
00050693
000c0593
000a8513
00068c13
2fc030ef
01012703
00050a93
000a0513
00070593
2e8030ef
00c12583
769020ef
00090593
2d8030ef
03812583
00050a13
000d8513
751020ef
000d0593
2c0030ef
00050d93
00098593
00048513
2b0030ef
00c12583
731020ef
00040593
2d5020ef
000d8593
298030ef
00050493
000c0593
00090513
2bd020ef
00050993
000a0593
000a8513
2ad020ef
00050713
000a0593
000a8513
00070a13
264030ef
00050a93
00090593
000c0513
254030ef
03c12583
00050c13
000b8513
6cd020ef
000d0593
271020ef
00048593
234030ef
00050d13
00040593
000d8513
224030ef
00050913
00098593
00040513
249020ef
67c030ef
00090593
00ab2023
000a0513
235020ef
668030ef
000a8593
00ab2223
00048513
221020ef
654030ef
000d0593
00ab2423
000c0513
20d020ef
640030ef
000d0593
00ab2623
000c0513
1c4030ef
62c030ef
00048593
00ab2823
000a8513
1b0030ef
618030ef
00090593
00ab2a23
000a0513
19c030ef
604030ef
00ab2c23
00040593
00098513
188030ef
5f0030ef
01412783
00ab2e23
000c8b13
d3979ae3
07c12083
07812403
07412483
07012903
06c12983
06812a03
06412a83
06012b03
05c12b83
05812c03
05412c83
05012d03
04c12d83
08010113
00008067
000217b7
a6c7a783
f8010113
06112e23
02f12623
000217b7
a747a783
06812c23
06912a23
02f12823
000217b7
a787a783
07212823
07312623
07412423
07512223
07612023
05712e23
05812c23
05912a23
05a12823
05b12623
02f12a23
00a12423
02b12c23
02c12e23
03812503
740010ef
01a00793
00a7cc63
03c12783
16078e63
03812503
728010ef
16a05863
00812683
000097b7
00008737
00e68733
00f687b3
24475703
8607a683
14e6f863
8567d403
8547c783
00001737
82170713
00e787b3
00812703
00479793
03f47413
00f707b3
68041e63
0047a483
03812903
00090513
76c010ef
000107b7
bff78793
64a7fc63
3ff57793
00179793
00f487b3
00001737
00e787b3
8017c583
00090513
8007c903
798010ef
00812703
000097b7
00f97993
00f707b3
8547c783
60079063
000087b7
25078793
00f707b3
00009a37
01470a33
856a5703
03812503
00098593
fc077713
00271713
00e784b3
65c010ef
00050813
0c041c63
02098063
fff98713
00100793
00e79733
00e55863
013797b3
fff78793
40f50533
00812603
00009737
00e605b3
8545c783
8565d683
00179793
00f607b3
00e787b3
85879603
03f6f713
00271713
00a60633
00e48733
00c72023
03812503
84c79c23
00168693
84d59b23
5e0010ef
01a00793
eaa7d2e3
00812683
000097b7
00008737
00e68733
00f687b3
24475703
8607a683
eae6ece3
07c12083
07812403
07412483
07012903
06c12983
06812a03
06412a83
06012b03
05c12b83
05812c03
05412c83
05012d03
04c12d83
00100513
08010113
00008067
856a5403
52091c63
03f47613
04060a63
00140693
000207b7
01069693
0106d693
9a078793
00c78633
00064703
00068413
03f6f613
00271713
00e48733
00168693
01069693
00072023
0106d693
fc061ce3
00812703
000097b7
00f707b3
84879b23
00812703
000097b7
00f707b3
8547c483
04000793
00049e63
000087b7
00f707b3
24b7c583
24a7c503
464030ef
00651793
daf440e3
00812683
00148793
00009737
00e68733
0ff7f793
00008437
84f70a23
84071b23
008684b3
2464ca03
d747eae3
24a4c583
24b4c503
424030ef
00050993
020508e3
00812783
2104ab03
35040413
00878933
00651b93
00000a93
f0090413
000b0493
0004d583
00042503
00440413
00248493
3e8030ef
fea42e23
fe8914e3
040a8a93
10090913
fd7a9ae3
00300793
7efa0463
00812783
00008437
25040493
009784b3
00000913
00878433
00048513
db0ff0ef
24b44583
24a44503
00190913
10048493
398030ef
fea942e3
24644703
00300793
7ef70e63
00812703
00008637
00c70bb3
24bbc783
2e078863
000217b7
a7c7a783
000096b7
00d70cb3
02f12423
000c8793
24abca03
000b8c93
00012823
00078b93
2c0a0263
01012783
00012623
0ff00993
00379a93
00279793
02f12223
000b8793
000c8b93
00078c93
00c12783
00000913
00379713
00279793
02f12023
000c8793
00e12a23
000b8c93
00078b93
0300006f
0ff00c93
01978123
24ad4c83
00140413
00800793
02f41863
00190913
000c8a13
000b0b93
000d0c93
20890c63
00391793
000c8d13
00f12223
00000413
000a0c93
000b8b13
850b5483
01412783
242d5c03
008484b3
00f484b3
fb84dae3
852b5783
240d5583
012787b3
01578a33
faba50e3
01012503
000c8593
280030ef
00c12783
00412703
00f507b3
00e405b3
00679793
00812703
00b787b3
00279793
00f707b3
246d4583
00008737
00f707b3
2507ad83
00300793
08f58263
080d8b93
000b8c93
000b8d93
000c0593
000a0513
22c030ef
00950533
864b2583
00151613
00a60633
00c585b3
0ff00793
0179c863
fffbc793
41f7d793
00fbf7b3
00f58023
864b2783
0ff00813
00c787b3
01b9c863
fffdc593
41f5d593
00bdf833
010780a3
864b2783
00c787b3
ed99cee3
fffcc613
41f65613
00ccfcb3
ed1ff06f
24bd4583
00090513
1dc030ef
02412783
000c8593
00f50cb3
00040513
1c8030ef
02012783
003c9c93
00f50533
00ac8cb3
000d8513
078030ef
00812783
002c9b93
00050c93
01778bb3
000087b7
01778bb3
750ba503
058030ef
02c12583
00a12e23
7f8020ef
000c8593
39c020ef
000217b7
a707a583
390020ef
7c5020ef
00050793
650ba503
00078b93
024030ef
03012583
00a12c23
7c4020ef
00050593
000c8513
331020ef
01c12883
03412583
00050d93
00088513
7a4020ef
00050593
000d8513
311020ef
000217b7
a707a583
338020ef
76d020ef
01812783
02812583
00050d93
00078513
774020ef
000c8593
318020ef
000217b7
a707a583
30c020ef
741020ef
00050c93
e89ff06f
00c12783
000d0b93
000b0c93
00178793
00f12623
d947c2e3
01012703
24bd4783
000d0c93
00170713
00e12823
000b0b93
d4f740e3
00812703
00009437
000087b7
00870433
86042503
00f707b3
2487d583
00150513
86a42023
00058663
0d0030ef
4e050863
00812703
000097b7
000086b7
00f707b3
84078a23
00d706b3
24a6c703
8507d583
2426d603
00371713
00b70733
01071713
01075713
84e79823
96c760e3
84079823
24b6c703
8527d683
00371713
00d70733
84e79923
945ff06f
00100713
38e78263
00812703
000087b7
75078793
00f707b3
9f9ff06f
00655793
01079793
0107d793
00179793
00f484b3
0014c583
03812503
0004c903
144010ef
9adff06f
0087a483
969ff06f
0f000793
34f90663
00495693
2e068063
000207b7
9a078793
03f47713
00e78733
00074703
00140613
01061613
00271713
00e48733
00100593
00072023
01065613
28b68263
03f67713
00e78733
00074583
00240713
01071713
00259593
00b485b3
00200893
0005a023
01075713
25168c63
03f77713
00e78733
00074583
00340713
01071713
00259593
00b485b3
00300893
0005a023
01075713
23168663
03f77593
00b785b3
0005c883
00170593
01059593
00289893
011488b3
00400313
0008a023
0105d593
20668063
03f5f593
00b785b3
0005c883
00270593
01059593
00289893
011488b3
00500313
0008a023
0105d593
1c668a63
03f5f593
00b785b3
0005c883
00370593
01059593
00289893
011488b3
00600313
0008a023
0105d593
1a668463
03f5f593
00b785b3
0005c883
00470593
01059593
00289893
011488b3
00700313
0008a023
0105d593
16668e63
03f5f593
00b785b3
0005c883
00570593
01059593
00289893
011488b3
00800313
0008a023
0105d593
14668863
03f5f593
00b785b3
0005c883
00670593
01059593
00289893
011488b3
00900313
0008a023
0105d593
12668263
03f5f593
00b785b3
0005c883
00770593
01059593
00289893
011488b3
00a00313
0008a023
0105d593
0e668c63
03f5f593
00b785b3
0005c883
00870593
01059593
00289893
011488b3
00b00313
0008a023
0105d593
0c668663
03f5f593
00b785b3
0005c883
00970593
01059593
00289893
011488b3
00c00313
0008a023
0105d593
0a668063
03f5f593
00b785b3
0005c883
00a70593
01059593
00289893
011488b3
00d00313
0008a023
0105d593
06668a63
03f5f593
00b785b3
0005c883
00b70593
01059593
00289893
011488b3
00e00313
0008a023
0105d593
04668463
03f5f593
00b785b3
0005c583
00c70713
01071713
00259593
00b485b3
01000893
0005a023
01075713
1b169a63
03f77713
00e78733
00074783
00279793
00f487b3
0007a023
00000793
00d05463
fff68793
00812703
00f60633
01061413
000097b7
01045413
00f707b3
84879b23
82098ce3
fff98713
00100793
00e79733
00e85863
013797b3
fff78793
40f80533
000207b7
03f47713
9a078793
00e787b3
0007c783
00140413
01041413
00279793
00f487b3
00a7a023
01045413
fdcff06f
00812703
000087b7
65078793
00f707b3
e78ff06f
000207b7
9a078793
00140613
03f47593
03f67713
00b785b3
0005c583
00240693
00e78733
00074703
03f6f693
00d786b3
0006c683
00259593
00b485b3
00271713
0005a023
00e48733
00072023
00269693
00340713
00d486b3
01061613
01071713
0006a023
01065613
01075713
01000693
cddff06f
00300793
86fa12e3
00812683
000087b7
00f68733
22072483
23072903
75078793
00f68433
08048a13
0004d583
f0042503
00290913
00440413
3b5020ef
ffe95583
00050793
ffc42503
eef42e23
00248493
39d020ef
fea42e23
fc9a18e3
fc099463
00812483
00008437
65040513
00a48533
d81fe0ef
75040513
00a48533
d75fe0ef
fe8ff06f
03812503
84042c23
84041e23
515000ef
b05ff06f
00f00693
e6dff06f
f7010113
00008737
08812423
08112623
08912223
09212023
07312e23
07412c23
07512a23
07612823
07712623
07812423
07912223
07a12023
05b12e23
00e50733
24070323
24071423
000057b7
08050023
00f507b3
20078623
000017b7
00f507b3
20078423
000067b7
10050123
00f507b3
200786a3
000027b7
00f507b3
200784a3
000077b7
18050223
00f507b3
20078723
000037b7
00f507b3
20078523
20050323
000047b7
200707a3
00f507b3
200785a3
000097b7
00f507b3
20070e23
22070623
22070e23
84078a23
84079b23
8407ac23
84079e23
8407a823
8607a023
86c7a223
0005c683
0ff00793
0015c603
00050413
0cf69663
0d800793
0cf61263
00100793
24f70623
ffff07b7
0ff78a93
ff0107b7
fff78b93
010007b7
00258493
fff78c13
000107b7
00001d37
bff78c93
00048913
00094683
0ff00713
00194783
10e69663
02078713
0ff77713
00f00693
0ae6fe63
0db00713
18e78463
0c000713
26e78863
0dd00713
0ee78c63
0c400713
38e78663
0da00713
7ce78263
0fe00713
12e78863
01078713
0ff77713
00d00693
12e6f063
0dc00713
10e78c63
02278713
0ff77713
00100693
10e6f463
34d78463
0ff00713
0ee79463
00390913
f79ff06f
000087b7
00f407b3
24078623
00000513
08c12083
08812403
08412483
08012903
07c12983
07812a03
07412a83
07012b03
06c12b83
06812c03
06412c83
06012d03
05c12d83
09010113
00008067
00294783
00394683
00490713
00879793
00d787b3
01079793
0107d793
ffe78613
00200693
00c70933
f0f6e0e3
00070913
00094683
0ff00713
00194783
eee68ee3
000087b7
00f407b3
24078623
00100513
f75ff06f
00294783
00394683
00494703
00594603
00879793
00d787b3
00871713
000086b7
00c70733
00d406b3
01079793
24e69423
0107d793
00400713
24e78263
000087b7
00f40433
24040623
00100513
f25ff06f
00294783
00394703
00200693
00879793
00e787b3
01079793
0107d793
00490713
f6f6f4e3
ffe78793
00f70933
e59ff06f
00294883
00394783
00490813
00889893
00f888b3
01089893
0108d893
ffe88893
09105263
00020e37
00100313
00084783
00180713
00c7f693
00f7f593
1c069463
0047d793
06078663
9a0e0613
00659513
04060f93
00b50f33
00064783
00074683
00174e83
00ff07b3
00179793
00869693
00f407b3
01d686b3
00160613
00d79023
00270713
fccf9ae3
08180813
f7f88893
00b507b3
00179793
00f407b3
08678023
f91046e3
f0089ce3
00080913
da9ff06f
9a0e0693
00659513
04068f13
00b50eb3
0006c783
00074603
00168693
00fe87b3
00179793
00f407b3
00c79023
00170713
fedf10e3
04180813
fbf88893
fa5ff06f
00494703
00800793
00294a03
00394d83
4cf71863
00594483
00694783
00008337
00849493
00f484b3
01049493
00640333
0104d493
24931023
00794503
00894703
00400793
00851513
00e50533
01051513
01055513
24a31123
00994983
00a90693
25330323
e6f984e3
48098c63
00199793
013787b3
00a78793
00f90933
00200e13
000088b7
00100813
00300e93
02c0006f
e3071ee3
e3039ce3
01178733
00659793
00b787b3
00179793
00f407b3
e2bee0e3
20f72023
45268863
0006c603
0016c703
00368693
00461793
fff60f13
00f407b3
00f77393
0fff7f13
011782b3
00839b13
00475f93
fff6c583
dfee62e3
20c2cf03
000f8713
016fefb3
dc0f1ae3
21028623
f90618e3
25f31523
f91ff06f
00690913
c55ff06f
00021537
83450513
1d5020ef
dadff06f
00290913
c3dff06f
00294783
00394683
00490713
00879793
00d787b3
01079793
0107d793
ffe78793
00f12a23
64f05c63
000047b7
20c78793
00f12e23
3ff00993
00812623
00074783
00c7f593
00f7f613
0047d693
34059a63
00c61793
00c787b3
36068663
01c12683
00d787b3
00c12683
00f68533
01a507b3
00100693
00d78023
00174583
00274483
00374f83
00474e03
009587b3
00574603
00674383
01f787b3
00774f03
01c787b3
00874303
00c787b3
00974683
007787b3
00a74283
01e787b3
00b74e83
00d74d83
00e74b03
006787b3
00c74883
00d787b3
00f74a03
005787b3
01d787b3
0156f6b3
015df833
00829293
008b1413
01074903
011787b3
0056e2b3
00849493
008866b3
0155f5b3
00839393
01567633
010a1813
0095e5b3
00766633
01b787b3
0176f6b3
0175f5b3
01767633
010e9e93
0106e6b3
010f9f93
010f1f13
0172f2b3
016787b3
01f5efb3
014787b3
01e665b3
0186f6b3
01d2e633
01891e93
012787b3
01d6e6b3
018e1e13
018ff833
01831313
0185f5b3
01889893
01867633
01c86833
0065e5b3
01166633
02d12a23
0ff7f693
03012423
02b12623
02c12823
00d12c23
0a200793
01170913
1ed7ee63
00250793
00f12823
000017b7
80278793
00900293
00100393
00000593
02810b13
01000a13
00f50433
007b07b3
fff7c303
0c030463
0ff3f613
ffa38f93
4079d4b3
41f9dfb3
407a0e33
00690333
00861f13
01861e93
01c597b3
00190913
fff94703
0cfcdc63
3ff7f793
01f7e833
06f84e63
40078693
00169693
00d506b3
0036fd93
40f808b3
120d9c63
0078bd93
120d9863
01577833
01e86833
01071d93
00188893
01787833
01b86833
0018dd93
01887833
002d9d93
01d86833
01b68db3
0106a023
00468693
fedd9ce3
ffe8f693
00f687b3
01168c63
00179793
00f507b3
01a787b3
80e78023
80c780a3
00158593
01059593
0105d593
f72310e3
00159593
01059593
00138393
01100793
0105d593
fff28293
f0f39ce3
01812783
01412703
01178793
0ff7f793
40f707b3
00f12a23
3cf05463
00090713
d61ff06f
005597b3
0097e833
0af9cc63
faf842e3
00179693
00d506b3
0036fd93
40f808b3
080d9063
0078bd93
060d9c63
01577833
01e86833
01071d93
00188893
01787833
01b86833
0018dd93
01887833
002d9d93
01d86833
01b68db3
0106a023
00468693
ffb69ce3
ffe8f693
00f687b3
f51682e3
00179793
00f507b3
00e78023
00c780a3
f31ff06f
00181793
008787b3
00e68023
00c680a3
00268693
fed79ae3
f15ff06f
00181793
01012803
010787b3
00e68023
00c680a3
00268693
fed79ae3
ef5ff06f
00c12403
000087b7
00f407b3
24078623
9adff06f
00021537
86050513
085020ef
9e1ff06f
00c12683
20878793
00f68533
c9dff06f
00068913
00008b37
01640b33
24ab4583
fff50513
008a1a13
00359593
288020ef
24bb4583
00050793
fff48513
00359593
00178493
270020ef
00150593
00048513
240020ef
ffed8793
014787b3
01079793
0107d793
00299713
24ab1223
ffa78793
41370733
80f700e3
965ff06f
000087b7
00f407b3
2467ce03
00294e83
00394603
00090493
8e0e0ce3
20078e23
00100713
00ee0e63
22078623
00200793
00fe0863
000087b7
00f407b3
22078e23
0044c683
00548793
08068a63
00169893
00588893
00004337
011488b3
000083b7
00100293
00300f93
20c30313
0540006f
20c74583
88059ee3
20570623
fff7c583
0045df13
00f5f813
00cf1513
00c5f493
00c81593
01e50533
010585b3
20850513
006585b3
00a40533
00b405b3
87efe2e3
860490e3
20a72223
20b72423
03178063
0007c583
00278793
00459713
00e40733
00770733
f8be7ee3
839ff06f
0007c583
0017c503
0027c703
820594e3
03f00593
82b510e3
80071ee3
008e9713
ffe60613
00e60633
00268713
01061693
0106d693
00171713
fee69e63
02810a13
000a0513
00008bb7
0037ca83
00478493
01740bb3
134000ef
24cbc783
0ff00b13
00700c93
0f800c13
02079a63
07c0006f
0c090663
03090793
0ff7f793
0afce863
0014ca83
00248493
000a0513
134000ef
02ac4c63
24cbc783
04078863
0004c903
00148993
fd6a86e3
000a8593
000a0513
0e8000ef
000a0513
00098493
00090a93
100000ef
fcac58e3
00000613
000a0593
00040513
941fe0ef
fa051ee3
000087b7
00f407b3
24078623
00100613
000a0593
00040513
921fe0ef
000087b7
00f407b3
04050a63
24c7c503
00154513
eacff06f
0009c903
00098493
03090793
0ff7f793
00090e63
f4fcfee3
00198993
ff6902e3
0d900793
faf914e3
fb1ff06f
0ff00593
000a0513
00248493
050000ef
fff4ca83
f39ff06f
24078623
00100513
e5cff06f
00070913
f2079063
000087b7
00f407b3
24c7c783
da079463
00100513
e3cff06f
00c12403
fe1ff06f
02051023
02050123
02052223
00008067
02054783
00f50733
00b70023
02452703
00178793
01f7f793
00870713
02f50023
02e52223
00008067
02452503
00008067
02154603
02254703
00800893
00260793
00160693
01f7f793
01f6f693
00d506b3
00f507b3
0006c803
0007c783
00c506b3
0006c683
40e888b3
00870313
4117d7b3
00e818b3
006696b3
0117e7b3
02452803
00b70733
00d7e7b3
01079793
40375693
01000893
40b888b3
00c686b3
0107d793
4117d7b3
01f6f693
00777713
40b80633
02d500a3
02e50123
02c52223
01079513
01055513
00008067
02154583
02254703
00258793
00158693
01f7f793
01f6f693
00d506b3
00f507b3
0007c783
0006c603
00b50533
00054683
00800593
40e585b3
40b7d533
00e617b3
00870713
00f56533
00e697b3
00f56533
01051513
01055513
00008067
02254783
02154603
02452683
00b787b3
4037d713
00c70733
01f77713
0077f793
40b686b3
02e500a3
02f50123
02d52223
00008067
02254703
02070663
02154783
02452683
00800613
40e60733
00178793
40e68733
01f7f793
02e52223
02050123
02f500a3
00008067
fb010113
05212023
0145d913
04912223
03312e23
03412c23
03512a23
03612823
00c59493
04112623
04812423
03712623
03812423
03912223
03a12023
01b12e23
7ff97913
00050993
00060b13
00068a93
00c4d493
01f5da13
0a090063
7ff00793
0ef90e63
01d55c93
00349493
009cecb3
008007b7
00fcecb3
00351413
c0190913
00000b93
014ad793
00ca9993
7ff7f793
00c9d993
01fada93
10078063
7ff00713
16e78063
00399993
01db5713
01376733
008009b7
013769b3
003b1813
c0178793
00000713
40f90933
002b9793
00e7e7b3
fff78793
00e00693
015a44b3
14f6ee63
000206b7
00279793
9e068693
00d787b3
0007a783
00078067
00a4ecb3
060c8e63
04048063
00048513
655010ef
ff550793
01c00713
02f74c63
01d00c93
ff850413
40fc8cb3
008494b3
0199dcb3
009cecb3
00899433
c0d00913
40a90933
f45ff06f
61d010ef
02050513
fc5ff06f
fd850c93
01999cb3
00000413
fddff06f
00a4ecb3
020c8463
00050413
00048c93
7ff00913
00300b93
f11ff06f
00000413
00000913
00100b93
f01ff06f
00000413
7ff00913
00200b93
ef1ff06f
0169e833
06080e63
04098063
00098513
5b5010ef
ff550713
01c00793
02e7ce63
01d00793
ff850813
40e787b3
010999b3
00fb57b3
0137e9b3
010b1833
c0d00793
40a787b3
ee5ff06f
000b0513
579010ef
02050513
fc1ff06f
fd850993
013b19b3
00000813
fd9ff06f
0169e833
02080263
000b0813
7ff00793
00300713
eb1ff06f
00000993
00000793
00100713
ea1ff06f
00000993
7ff00793
00200713
e91ff06f
0199e663
453c9a63
45046863
01fc9713
00145793
01f41d93
001cdc93
00f76433
01885a93
00899b93
017aeab3
010bdb93
000b8593
010a9c13
000c8513
00881b13
010c5c13
3c5010ef
00050593
00050d13
000c0513
389010ef
00050993
000b8593
000c8513
3ed010ef
01051513
01045713
00a76733
000d0a13
01377e63
01570733
fffd0a13
01576863
01377663
ffed0a13
01570733
413709b3
000b8593
00098513
369010ef
00050593
00050d13
000c0513
32d010ef
00050c93
000b8593
00098513
391010ef
01041413
01051513
01045413
00a46433
000d0793
01947e63
01540433
fffd0793
01546863
01947663
ffed0793
01540433
010a1713
00010337
00f76733
41940433
fff30c93
019777b3
019b7cb3
01075e13
010b5d13
00078513
000c8593
2bd010ef
00050813
000d0593
00078513
2ad010ef
00050793
000c8593
000e0513
29d010ef
00050893
000d0593
000e0513
28d010ef
01085a13
011787b3
00fa0a33
00050693
011a7463
006506b3
010a5793
00d787b3
000106b7
fff68693
00da7a33
010a1a13
00d87833
010a0a33
00f46863
00070993
04f41463
054df263
016d8db3
016db6b3
015686b3
00d40433
fff70993
008ae663
028a9463
036de263
00f46663
00879e63
014dfc63
016d8db3
ffe70993
016db733
01570733
00e40433
414d8a33
40f40433
014db7b3
40f40433
fff00813
1a8a8263
000b8593
00040513
20d010ef
00050593
00a12623
000c0513
1d1010ef
00a12423
000b8593
00040513
235010ef
00c12683
00812783
01051513
010a5713
00a76733
00068d93
00f77e63
01570733
fff68d93
01576863
00f77663
ffe68d93
01570733
40f70433
000b8593
00040513
1a9010ef
00050593
00a12423
000c0513
16d010ef
00050c13
000b8593
00040513
1d1010ef
00812783
010a1713
01051513
01075713
00a76733
00078693
01877e63
01570733
fff78693
01576863
01877663
ffe78693
01570733
010d9793
00d7e7b3
01079813
01085813
41870733
0107de13
00080513
000c8593
105010ef
00050893
000d0593
00080513
0f5010ef
00050813
000c8593
000e0513
0e5010ef
00050313
000d0593
000e0513
0d5010ef
0108d693
00680833
010686b3
00050593
0066f663
00010637
00c505b3
0106d613
00b60633
000105b7
fff58593
00b6f6b3
01069693
00b8f8b3
011686b3
00c76863
24c71a63
00078813
04068063
00ea8733
fff78813
03576463
00c76663
22c71a63
02db7063
ffe78813
001b1793
0167bb33
015b0b33
01670733
00078b13
00c71463
00db0463
00186813
3ff90793
12f05063
00787713
02070063
00f87713
00400693
00d70a63
00480713
01073833
010989b3
00070813
01000737
00e9f733
00070a63
ff0007b7
fff78793
00f9f9b3
40090793
7fe00713
0af74663
00385813
01d99713
01076733
0039d593
7ff006b7
01479793
00c59593
04c12083
04812403
00d7f7b3
00c5d593
00b7e7b3
01f49493
0097e6b3
04012903
04412483
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
00070513
00068593
05010113
00008067
fff90913
00000d93
bc1ff06f
000a0493
000c8993
00040813
000b8713
00300793
10f70063
00100793
0ef70663
00200793
f0f716e3
00000593
00000713
7ff00793
f5dff06f
000a8493
fd5ff06f
000809b7
00000813
00000493
00300713
fc1ff06f
00100593
40f585b3
03800713
0ab74463
01f00713
06b74663
41e90913
012997b3
00b85733
01281933
00e7e7b3
01203933
0127e7b3
00b9d5b3
0077f713
02070063
00f7f713
00400693
00d70a63
00478713
00f737b3
00f585b3
00070793
00800737
00e5f733
06071863
01d59713
0037d793
00f76733
0035d593
00000793
ec1ff06f
fe100713
40f707b3
02000693
00f9d7b3
00000713
00d58663
43e90713
00e99733
01076733
00e03733
00e7e7b3
00000593
f89ff06f
00000593
00000713
fbdff06f
000805b7
00000713
7ff00793
00000493
e6dff06f
00000593
00000713
00100793
e5dff06f
00080793
00078813
dedff06f
fd010113
01312e23
0145d993
02812423
02912223
01412c23
01512a23
01712623
00c59493
02112623
03212023
01612823
7ff9f993
00050413
00060b93
00068a13
00c4d493
01f5da93
3c098863
7ff00793
42f98663
00349493
01d55793
0097e7b3
008004b7
0097e4b3
00351913
c0198993
00000b13
014a5713
00ca1413
7ff77713
00c45413
01fa5a13
42070663
7ff00793
48f70663
00341413
01dbd793
0087e7b3
00800437
0087e433
c0170713
003b9793
00000613
00e989b3
002b1713
00c76733
00a00693
014ac833
00198893
4ce6c863
00200693
48e6c063
fff70713
00100693
48e6fc63
00010a37
fffa0393
0107d293
00797e33
0077f7b3
01095f93
000e0513
00078593
530010ef
00050e93
00028593
000e0513
520010ef
00050713
00078593
000f8513
510010ef
00050913
00028593
000f8513
500010ef
010ed313
01270733
00e30333
00050f13
01237463
01450f33
01035913
00737333
007efeb3
01031313
007473b3
01d30333
01045a13
000e0513
00038593
4c0010ef
00050e93
000a0593
000e0513
4b0010ef
00050e13
00038593
000f8513
4a0010ef
00050413
000a0593
000f8513
490010ef
010ed713
008e0e33
01c70733
00050693
00877663
00010637
00c506b3
00010b37
fffb0e13
01075f93
01c77733
01071713
01cefeb3
01d70eb3
01c4fe33
00df8fb3
01d90933
0104da93
000e0513
00078593
43c010ef
00050413
00028593
000e0513
42c010ef
00050493
00078593
000a8513
41c010ef
00050b93
00028593
000a8513
40c010ef
01045793
017484b3
009787b3
00050713
0177f463
01650733
000104b7
fff48693
0107d293
00e282b3
00d7f733
00d47433
01071713
00870733
000e0513
00038593
3c8010ef
00050413
000a0593
000e0513
3b8010ef
00050e13
00038593
000a8513
3a8010ef
00050393
000a0593
000a8513
398010ef
01045793
007e0e33
01c78e33
00050593
007e7463
009505b3
000106b7
fff68693
00de77b3
00d47433
01079793
012f0f33
008787b3
01df3eb3
01f787b3
01d78533
00ef0f33
00ef3733
005506b3
00e68633
01f7b433
01d53533
010e5793
00e63733
00a46433
0056b6b3
00f40433
00e6e6b3
00d40433
00b40433
01765793
00941413
00f46433
009f1793
0067e7b3
00f037b3
017f5f13
00961713
01e7e7b3
00e7e7b3
01000737
00e47733
28070663
0017d713
0017f793
00f76733
01f41793
00f767b3
00145413
3ff88693
26d05a63
0077f713
02070063
00f7f713
00400613
00c70a63
00478713
00f737b3
00f40433
00070793
01000737
00e47733
00070a63
ff000737
fff70713
00e47433
40088693
7fe00713
2ed74e63
01d41713
0037d793
00f76733
00345413
7ff007b7
01469693
00c41413
00f6f6b3
00c45413
02c12083
0086e6b3
02812403
01f81813
0106e7b3
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00070513
00078593
03010113
00008067
00a4e933
06090c63
04048063
00048513
354010ef
ff550713
01c00793
02e7cc63
01d00793
ff850913
40e787b3
012494b3
00f457b3
0097e4b3
01241933
c0d00993
40a989b3
c15ff06f
31c010ef
02050513
fc5ff06f
fd850493
009414b3
00000913
fddff06f
00a4e933
02090263
00050913
7ff00993
00300b13
be5ff06f
00000493
00000993
00100b13
bd5ff06f
00000493
7ff00993
00200b13
bc5ff06f
017467b3
06078e63
04040063
00040513
2b8010ef
ff550693
01c00793
02d7ce63
01d00713
ff850793
40d70733
00f41433
00ebd733
00876433
00fb97b3
c0d00713
40a70733
bb9ff06f
000b8513
27c010ef
02050513
fc1ff06f
fd850413
008b9433
00000793
fd9ff06f
017467b3
02078263
000b8793
7ff00713
00300613
b85ff06f
00000413
00000713
00100613
b75ff06f
00000413
7ff00713
00200613
b65ff06f
00100693
00e696b3
5306f713
04071863
2406f593
12059463
0886f693
b6068ae3
000a0813
00200713
12e60863
00300713
10e60e63
00100713
dce61ce3
00000413
00000713
0bc0006f
00f00693
02d70063
00b00693
fcd706e3
000a8813
00048413
00090793
000b0613
fbdff06f
00080437
00000793
00000813
00300613
fb1ff06f
00098893
d8dff06f
00100613
40d60633
03800713
fac744e3
01f00713
06c74663
41e88893
01141733
00c7d6b3
011798b3
00d76733
011038b3
011767b3
00c45433
0077f713
02070063
00f7f713
00400693
00d70a63
00478713
00f737b3
00f40433
00070793
00800737
00e47733
06071e63
01d41713
0037d793
00f76733
00345413
00000693
d6dff06f
fe100713
40d70733
02000593
00e45733
00000693
00b60663
43e88893
011416b3
00f6e6b3
00d036b3
00d767b3
00000413
f89ff06f
00080437
7ff00693
00000813
d29ff06f
00080437
00000713
fedff06f
00000413
00000713
7ff00693
d0dff06f
00000413
00000713
00100693
cfdff06f
fe010113
00112e23
00812c23
00912a23
01212823
01312623
01412423
00b567b3
16078e63
00050413
00058913
00058493
08058463
00058513
078010ef
00050993
43e00a13
413a0a33
43300793
0947c463
00b00713
00040793
02e98463
02a00713
07374263
02b00493
ff598713
413484b3
009454b3
00e91933
0124e4b3
00e417b3
01c12083
01812403
00c49593
014a1a13
00c5d593
00ba6733
01412483
01012903
00c12983
00812a03
00078513
00070593
02010113
00008067
7f9000ef
02050993
f81ff06f
fd598593
00b414b3
00000793
fb1ff06f
43600793
0347dc63
03898613
00040513
00090593
791000ef
00b56533
00800613
00a034b3
00090593
00040513
41360633
73d000ef
00a4e433
00058913
00800713
00040793
03375063
02800713
ff898693
41370733
00d91933
00e45733
01276933
00d417b3
ff800737
fff70713
00e975b3
0077f713
02070063
00f7f713
00400693
00d70a63
00478713
00f737b3
00f585b3
00070793
00800737
00e5f733
00070c63
ff800737
fff70713
43f00a13
00e5f5b3
413a0a33
0037d793
01d59713
00f767b3
0035d493
ee9ff06f
00000493
00000793
00000a13
ed9ff06f
00800737
ff010113
fff70713
00a777b3
00812423
00912223
01755413
01f55493
0175d513
00b77733
0ff47413
0ff57513
00112623
01212023
01f5d593
00379793
00371713
40a406b3
18b49663
0ad05863
04051063
02070063
fff40693
00069863
00e787b3
00100413
0600006f
0ff00613
02c41863
0077f713
34070a63
00f7f713
00400693
34d70463
00478793
3400006f
0ff00613
fec400e3
04000637
00c76733
01b00593
00100613
00d5ce63
02000613
00d755b3
40d606b3
00d71733
00e03733
00e5e633
00c787b3
04000737
00e7f733
fa0702e3
00140413
0ff00713
2ee40663
7e000737
0017f693
fff70713
0017d793
00e7f7b3
00d7e7b3
f7dff06f
06068663
408506b3
02041063
2a078663
fff68613
f40608e3
0ff00593
02b69063
00070793
2100006f
0ff00613
fec50ae3
04000637
00c7e7b3
00068613
01b00593
00100693
00c5ce63
02000693
40c686b3
00c7d5b3
00d797b3
00f037b3
00f5e6b3
00e687b3
00050413
f65ff06f
00140693
0fe6f613
04061663
02041863
24078263
ee070ce3
00e787b3
04000737
00e7f733
ee0704e3
fc000737
fff70713
00e7f7b3
00100413
ed5ff06f
f6078ce3
18070463
00000493
020007b7
0ff00413
2140006f
0ff00613
20c68263
00e78733
00175793
00068413
ea5ff06f
06d05e63
06051263
e8070ce3
fff40693
00069863
40e787b3
00100413
0340006f
0ff00613
e6c40ee3
01b00593
00100613
00d5ce63
02000613
00d755b3
40d606b3
00d71733
00e03733
00e5e633
40c787b3
04000937
0127f733
e40704e3
fff90913
0127f933
1180006f
0ff00613
e2c40ae3
04000637
00c76733
fb1ff06f
08068063
408506b3
02041863
1e078263
fff68613
00061863
40f707b3
00058493
f7dff06f
0ff00813
03069263
00070793
0ff00413
06c0006f
0ff00613
fec508e3
04000637
00c7e7b3
00068613
01b00813
00100693
00c84e63
02000693
40c686b3
00c7d833
00d797b3
00f037b3
00f866b3
40d707b3
00050413
00058493
f59ff06f
00140693
0fe6f693
06069063
04041263
00079c63
00000493
0e070263
00070793
00058493
d81ff06f
d6070ee3
40e786b3
04000637
00c6f633
40f707b3
fe0612e3
00000793
08068263
00068793
d59ff06f
e80794e3
e80704e3
00070793
00058493
0ff00413
d41ff06f
40e78933
040006b7
00d976b3
04068463
40f70933
00058493
00090513
3b1000ef
ffb50513
00a91933
04854063
40850533
00150513
02000713
40a70733
00a957b3
00e91933
01203933
0127e7b3
00000413
cedff06f
fc0912e3
00000793
00000413
00000493
0300006f
fc0007b7
fff78793
40a40433
00f977b3
cc5ff06f
00070793
e15ff06f
00070793
cb5ff06f
0ff00413
00000793
04000737
00e7f733
00070e63
00140413
0ff00713
06e40663
fc000737
fff70713
00e7f7b3
0ff00713
0037d793
00e41863
00078663
004007b7
00000493
01741413
7f800737
00979793
00e47433
0097d793
00f46433
01f49513
00c12083
00a46533
00812403
00412483
00012903
01010113
00008067
00070793
00068413
ea9ff06f
00000793
fa1ff06f
fe010113
01212823
01755913
00912a23
01312623
01512223
00951493
00112e23
00812c23
01412423
0ff97913
00058a93
0094d493
01f55993
1c090263
0ff00793
1cf90e63
00349493
040007b7
00f4e4b3
f8190913
00000a13
017ad793
009a9413
0ff7f793
00945413
01fada93
1c078863
0ff00713
1ee78463
00341413
04000737
00e46433
f8178793
00000693
00f90933
002a1793
00d7e7b3
00a00713
0159c833
00190893
22f74463
00200713
1cf74863
fff78793
00100713
1ef77463
00010eb7
fffe8313
0104df93
01045f13
0064f4b3
00647433
00048513
00040593
08d000ef
00050713
000f0593
00048513
07d000ef
00050793
00040593
000f8513
06d000ef
00050e13
000f0593
000f8513
05d000ef
01075413
01c787b3
00f40433
00050693
01c47463
01d506b3
006477b3
00677733
01079793
00e787b3
00679713
01045413
00e03733
01a7d793
00d40433
00f767b3
00641413
00f46433
080007b7
00f477b3
18078e63
00145793
00147413
0087e433
07f88713
18e05863
00747793
00078a63
00f47793
00400693
00d78463
00440413
080007b7
00f477b3
00078a63
f80007b7
fff78793
00f47433
08088713
0fe00793
1ae7ce63
00345793
01c12083
01812403
01771713
7f8006b7
00979793
00d77733
0097d793
00f76733
01f81513
01412483
01012903
00c12983
00812a03
00412a83
00a76533
02010113
00008067
02048a63
00048513
0ad000ef
ffb50793
f8a00913
00f494b3
40a90933
e3dff06f
0ff00913
00200a13
e2048ae3
00300a13
e2dff06f
00000913
00100a13
e21ff06f
02040a63
00040513
06d000ef
ffb50793
00f41433
f8a00793
40a787b3
e31ff06f
0ff00793
00200693
e20404e3
00300693
e21ff06f
00000793
00100693
e15ff06f
00100713
00f717b3
5307f713
04071c63
2407f713
0c071663
0887f793
e20782e3
000a8813
00200613
00000793
0ff00713
f0c686e3
00300793
0af68463
00100793
eaf69ae3
00000793
00000713
ef1ff06f
00f00713
00e78e63
00b00713
fce782e3
00098813
00048413
000a0693
fb9ff06f
00400437
00000813
00300693
fb9ff06f
00090893
e71ff06f
00100793
40e787b3
01b00713
faf748e3
09e88893
00f457b3
01141433
00803433
0087e7b3
0077f713
00070a63
00f7f713
00400693
00d70463
00478793
04000737
00e7f733
0037d793
e60706e3
00000793
00100713
e61ff06f
004007b7
0ff00713
00000813
e51ff06f
00000793
0ff00713
e45ff06f
00800737
ff010113
fff70713
0175d613
00a777b3
00812423
00b77733
00912223
01755413
00112623
01212023
0ff67613
0ff00693
0ff47413
01f55493
00379793
01f5d593
00371713
00d61463
00071463
0015c593
40c406b3
18959a63
0ad05063
02061663
18070063
fff68613
00061863
00e787b3
00100413
0500006f
0ff00593
02b69063
0ff00413
1180006f
0ff00613
10c40863
04000637
00c76733
00068613
01b00593
00100693
00c5ce63
02000693
40c686b3
00c755b3
00d71733
00e03733
00e5e6b3
00d787b3
04000737
00e7f733
0c070863
00140413
0ff00713
30e40263
7e000737
0017f693
fff70713
0017d793
00e7f7b3
00d7e7b3
0a80006f
06068663
408606b3
02041063
2c078263
fff68593
f60580e3
0ff00513
02a69063
00070793
f65ff06f
0ff00593
feb60ae3
040005b7
00b7e7b3
00068593
01b00513
00100693
00b54e63
02000693
40b686b3
00b7d533
00d797b3
00f037b3
00f566b3
00e687b3
00060413
f65ff06f
00140693
0fe6f613
06061263
04041463
24078e63
02070263
00e787b3
04000737
00e7f733
00070a63
fc000737
fff70713
00e7f7b3
00100413
0077f713
24070063
00f7f713
00400693
22d70a63
00478793
22c0006f
f60780e3
ec0702e3
00000493
020007b7
0ff00413
2140006f
0ff00613
20c68263
00e78733
00175793
00068413
fb9ff06f
08d05063
06061263
fe0708e3
fff68613
00061863
40e787b3
00100413
0340006f
0ff00593
e6b68ae3
01b00593
00100693
00c5ce63
02000693
40c686b3
00c755b3
00d71733
00e03733
00e5e6b3
40d787b3
04000937
0127f733
f4070ee3
fff90913
0127f933
1180006f
0ff00613
f4c404e3
04000637
00c76733
00068613
fadff06f
08068063
408606b3
02041863
1e078063
fff68513
00051863
40f707b3
00058493
f79ff06f
0ff00813
03069263
00070793
0ff00413
06c0006f
0ff00513
fea608e3
04000537
00a7e7b3
00068513
01b00813
00100693
00a84e63
02000693
40a686b3
00a7d833
00d797b3
00f037b3
00f866b3
40d707b3
00060413
00058493
f55ff06f
00140693
0fe6f693
04069e63
04041263
00079c63
00000493
0e070063
00070793
00058493
e91ff06f
e80706e3
40e786b3
04000637
00c6f633
40f707b3
fe0612e3
00000793
08068063
00068793
e69ff06f
e80792e3
e80702e3
00070793
00058493
d39ff06f
40e78933
040006b7
00d976b3
04068463
40f70933
00058493
00090513
3cc000ef
ffb50513
00a91933
04854063
40850533
00150513
02000713
40a70733
00a957b3
00e91933
01203933
0127e7b3
00000413
e01ff06f
fc0912e3
00000793
00000413
00000493
0300006f
fc0007b7
fff78793
40a40433
00f977b3
dd9ff06f
00070793
e15ff06f
00070793
dc9ff06f
0ff00413
00000793
04000737
00e7f733
00070e63
00140413
0ff00713
06e40663
fc000737
fff70713
00e7f7b3
0ff00713
0037d793
00e41863
00078663
004007b7
00000493
01741413
7f800737
00979793
00e47433
0097d793
00f46433
01f49513
00c12083
00a46533
00812403
00412483
00012903
01010113
00008067
00070793
00068413
eadff06f
00000793
fa1ff06f
00800637
01755713
fff60793
0ff77713
07e00593
00a7f7b3
01f55693
04e5d663
09d00593
00e5da63
80000537
fff54513
00a68533
00008067
00c7e533
09500793
00e7dc63
f6a70713
00e51533
02068063
40a00533
00008067
09600793
40e787b3
00f55533
fe9ff06f
00000513
00008067
0e050863
41f55793
ff010113
00812423
00a7c433
40f40433
00912223
01f55493
00040513
00112623
234000ef
09e00713
40a70733
09600793
02e7cc63
ff850513
00a417b3
00c12083
00812403
00979793
01771713
0097d793
01f49513
00f76733
00412483
00a76533
01010113
00008067
09900793
02e7d063
00500793
40a787b3
01b50693
00f457b3
00d41433
00803433
0087e433
00500793
00a7d663
ffb50793
00f41433
fc0007b7
fff78793
00747693
00f477b3
00068a63
00f47413
00400693
00d40463
00478793
040006b7
00d7f6b3
00068c63
fc000737
fff70713
00e7f7b3
09f00713
40a70733
0037d793
f59ff06f
00000793
00000713
00979793
0097d793
01771713
00f76733
01f51513
00a76533
00008067
00050613
00000513
0015f693
00068463
00c50533
0015d593
00161613
fe0596e3
00008067
06054063
0605c663
00058613
00050593
fff00513
02060c63
00100693
00b67a63
00c05863
00161613
00169693
feb66ae3
00000513
00c5e663
40c585b3
00d56533
0016d693
00165613
fe0696e3
00008067
00008293
fb5ff0ef
00058513
00028067
40a00533
00b04863
40b005b3
f9dff06f
40b005b3
00008293
f91ff0ef
40a00533
00028067
00008293
0005ca63
00054c63
f79ff0ef
00058513
00028067
40b005b3
fe0558e3
40a00533
f61ff0ef
40b00533
00028067
02060063
02000793
40c787b3
00f04c63
fe060613
00c5d533
00000713
00070593
00008067
00c5d733
00c55533
00f595b3
00b56533
fe9ff06f
02060063
02000793
40c787b3
00f04c63
fe060613
00c515b3
00000713
00070513
00008067
00c51733
00c595b3
00f55533
00a5e5b3
fe9ff06f
000107b7
02f57a63
10053793
0017c793
00379793
00020737
02000693
40f686b3
00f55533
a1c70793
00a787b3
0007c503
40a68533
00008067
01000737
01000793
fce56ae3
01800793
fcdff06f
ff010113
00000593
00812423
00112623
00050413
118030ef
000217b7
a2c7a503
03c52783
00078463
000780e7
00040513
4350f0ef
ff010113
00812423
01212023
00000793
00000913
40f90933
00112623
00912223
40295913
02090063
00000413
00000493
00042783
00148493
00440413
000780e7
fe9918e3
00000793
00000913
40f90933
40295913
02090063
00000413
00000493
00042783
00148493
00440413
000780e7
fe9918e3
00c12083
00812403
00412483
00012903
01010113
00008067
00f00313
00050713
02c37e63
00f77793
0a079063
08059263
ff067693
00f67613
00e686b3
00b72023
00b72223
00b72423
00b72623
01070713
fed766e3
00061463
00008067
40c306b3
00269693
00000297
005686b3
00c68067
00b70723
00b706a3
00b70623
00b705a3
00b70523
00b704a3
00b70423
00b703a3
00b70323
00b702a3
00b70223
00b701a3
00b70123
00b700a3
00b70023
00008067
0ff5f593
00859693
00d5e5b3
01059693
00d5e5b3
f6dff06f
00279693
00000297
005686b3
00008293
fa0680e7
00028093
ff078793
40f70733
00f60633
f6c378e3
f3dff06f
fc010113
02c12423
02d12623
02e12823
02f12a23
03012c23
03112e23
00058613
00852583
02810693
00112e23
00d12623
328000ef
01c12083
04010113
00008067
04007337
67432303
fc010113
02c12423
02d12623
02b12223
02e12823
02f12a23
03012c23
03112e23
00832583
02410693
00050613
00030513
00112e23
00d12623
2d8000ef
01c12083
04010113
00008067
00852603
01c0006f
040077b7
6747a783
00050593
0087a603
00078513
0040006f
fe010113
01212c23
00112e23
00050913
00050663
03852783
04078663
00862783
fff78793
00f62423
0007dc63
01862703
04e7c663
0ff5f793
00a00713
04e78063
00062783
0ff5f513
00178713
00e62023
00b78023
01c12083
01812903
02010113
00008067
00c12623
00b12423
644030ef
00c12603
00812583
fa5ff06f
01c12083
00090513
01812903
02010113
3490206f
ff010113
040077b7
01212023
6747a903
00812423
00912223
00112623
00050493
00058413
00090663
03892783
04078a63
00842783
fff78793
00f42423
0007dc63
01842703
04e7c463
0ff4f793
00a00713
02e78e63
00042783
0ff4f513
00178713
00e42023
00978023
00c12083
00812403
00412483
00012903
01010113
00008067
00090513
59c030ef
fa9ff06f
00040613
00812403
00c12083
00048593
00090513
00412483
00012903
01010113
2990206f
fc010113
02812c23
00050413
00058513
02912a23
02112e23
00058493
0c0000ef
000207b7
74c78793
02f12423
00100793
02f12623
03842703
02010793
00150693
00f12a23
00200793
02912023
02a12223
00d12e23
00f12c23
00842583
04070e63
00c59783
01279713
02074263
0645a703
000026b7
00d7e7b3
ffffe6b7
fff68693
00d77733
00f59623
06e5a223
01410613
00040513
1cd030ef
03c12083
03812403
00a03533
40a00533
03412483
00a56513
04010113
00008067
00040513
00b12623
4b0030ef
00c12583
f99ff06f
040077b7
00050593
6747a503
f29ff06f
00357793
00050713
04079c63
7f7f86b7
f7f68693
fff00593
00072603
00470713
00d677b3
00d787b3
00c7e7b3
00d7e7b3
feb784e3
ffc74683
40a707b3
04068463
ffd74683
02068c63
ffe74503
00a03533
00f50533
ffe50513
00008067
fa0688e3
00074783
00170713
00377693
fe0798e3
40a70733
fff70513
00008067
ffd78513
00008067
ffc78513
00008067
e1010113
1e112623
1f212023
1d812423
1da12023
00058c13
00060913
00d12a23
1e812423
1e912223
1d312e23
1d412c23
1d512a23
1d612823
1d712623
1d912223
1bb12e23
00050d13
251060ef
00052783
00078513
02f12823
f1dff0ef
02a12623
0e012823
0e012a23
0e012c23
0e012e23
000d0663
038d2783
70078863
00cc1683
00002637
01069793
0107d793
00c7f5b3
02059863
064c2583
00c6e7b3
01079793
ffffe6b7
4107d793
fff68693
00d5f6b3
00fc1623
01079793
06dc2223
0107d793
0087f693
2e068663
010c2683
2e068263
01a7f793
00a00693
2ed78e63
10c10793
00078893
0ef12223
000207b7
c2078793
00f12c23
000207b7
e3478793
00090b13
00f12423
000b4783
0e012623
0e012423
02012023
02012a23
02012c23
02012e23
04012223
04012423
00012623
00088c93
22078263
000b0413
02500713
30e78463
00144783
00140413
fe079ae3
416404b3
21640263
0ec12703
0e812783
016ca023
00970733
00178793
009ca223
0ee12623
0ef12423
00700713
008c8c93
2cf74c63
00c12703
00044783
00970733
00e12623
1c078263
fff00313
00144483
0c0103a3
00140413
00000993
00000a13
05a00913
00900a93
02a00b93
00030d93
00140413
fe048793
04f96463
01812703
00279793
00e787b3
0007a783
00078067
00000993
fd048693
00044483
00299793
013787b3
00179793
00f689b3
fd048693
00140413
fedaf2e3
fe048793
fcf970e3
14048463
14910623
0c0103a3
00100a93
00100b93
14c10b13
00012823
00000313
02012423
02012223
00012e23
002a7f93
000f8463
002a8a93
084a7913
0ec12783
00091663
415986b3
44d04ee3
0c714703
02070a63
0e812703
0c710693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
2ee6ca63
020f8a63
0e812703
0c810693
00dca023
00278793
00200693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
52e6c0e3
08000713
22e900e3
41730db3
31b040e3
100a7713
0c071ee3
0e812703
017787b3
016ca023
00170713
017ca223
0ef12623
0ee12423
00700693
3ae6ce63
008c8c93
004a7a13
000a0663
415984b3
3c904463
0159d463
000a8993
00c12703
01370733
00e12623
360790e3
01012783
0e012423
00078863
01012583
000d0513
2a4030ef
10c10c93
00040b13
000b4783
de0792e3
0ec12783
00078463
2ed0106f
00cc5783
0407f793
00078463
2240206f
1ec12083
1e812403
00c12503
1e412483
1e012903
1dc12983
1d812a03
1d412a83
1d012b03
1cc12b83
1c812c03
1c412c83
1c012d03
1bc12d83
1f010113
00008067
000c0593
000d0513
714020ef
00050463
1d00206f
00cc5783
00a00693
01a7f793
d0d796e3
00ec1783
d007c2e3
01412683
00090613
000c0593
000d0513
480020ef
00a12623
f7dff06f
000d0513
69c060ef
00452783
00078513
04f12423
b69ff0ef
00050793
000d0513
00078493
04f12223
678060ef
00852783
02f12e23
720492e3
00044483
d89ff06f
00044483
020a6a13
d7dff06f
416404b3
d16416e3
00044783
d41ff06f
0e410613
000c0593
000d0513
4150b0ef
ee051ee3
10c10c93
d15ff06f
008a7793
000d8313
70079ee3
01412783
0b010513
01b12823
00778793
ff87f793
0047a603
0007a583
00878793
00f12a23
5e1120ef
0b012603
0b412683
0b812703
0bc12783
01012303
0f010513
00612823
0ef12e23
0ec12823
0ed12a23
0ee12c23
548060ef
0ca12623
00200793
01012303
00f51463
2900106f
00100793
00f51463
3e00106f
06100793
00f49463
7650106f
04100793
00f49463
1850106f
fdf4f713
fff00793
02e12423
00f31463
19c0206f
04700793
00f71463
1800206f
0fc12d83
05412023
0f012e03
0f412e83
0f812f03
100a6793
000dd463
6b90106f
04012c23
00078a13
00012823
fbf48793
02500713
00f77463
5fc0106f
00020737
00279793
d8c70713
00e787b3
0007a783
00078067
0e410613
000c0593
000d0513
04612623
05f12023
2e10b0ef
100512e3
0ec12783
04c12303
04012f83
10c10c93
ce5ff06f
0e812483
02012683
00100713
016ca023
00178793
00148493
008c8d93
3ad75ae3
00100713
00eca223
0ef12623
0e912423
00700713
769740e3
02c12703
03012683
00148493
00e787b3
00eda223
00dda023
0ef12623
0e912423
00700713
008d8d93
74974ce3
0f012703
0a010593
0b010513
0ae12823
0f412703
00f12e23
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
5950f0ef
02012783
fff78913
01c12783
360500e3
001b0813
00148493
012787b3
010da023
012da223
0ef12623
0e912423
00700713
008d8d93
30974ae3
03812683
0d410713
00148493
00f687b3
00eda023
00dda223
0ef12623
0e912423
00700713
008d8c93
c49758e3
0e410613
000c0593
000d0513
1b10b0ef
7c051a63
0ec12783
10c10c93
c31ff06f
01000693
0e812703
0096c463
6710106f
000206b7
e2468d93
01000913
00700a13
00c0006f
ff048493
04995663
01078793
00170713
01bca023
012ca223
0ef12623
0ee12423
008c8c93
fcea5ee3
0e410613
000c0593
000d0513
1450b0ef
76051463
ff048493
0ec12783
0e812703
10c10c93
fa994ee3
009787b3
00170713
01bca023
009ca223
0ef12623
0ee12423
00700693
bae6d6e3
0e410613
000c0593
000d0513
0fd0b0ef
72051063
0ec12783
b91ff06f
000d0513
47d020ef
8edff06f
01412703
0c0103a3
00100a93
00072783
00470713
00e12a23
14f10623
00100b93
14c10b13
a6dff06f
01412783
0c0103a3
0007ab03
00478913
4c0b00e3
fff00793
00fd9463
04c0106f
000d8613
00000593
000b0513
01b12a23
661060ef
00a12823
01412303
00051463
4ad0106f
01012783
41678bb3
0c714783
fffbca93
41fada93
01212a23
00012823
02012423
02012223
00012e23
015bfab3
00000313
a00784e3
001a8a93
a01ff06f
01412783
0007a983
00478793
2a09d8e3
413009b3
00f12a23
00044483
004a6a13
961ff06f
01412683
020a7793
00468713
300794e3
010a7793
780790e3
040a7793
00078463
5740106f
200a7a13
760a06e3
01412783
00e12a23
00c12703
0007a783
00040b13
00e78023
aa9ff06f
00044483
06c00793
38f48ee3
010a6a13
905ff06f
01412703
ffff87b7
8307c793
0cf11423
00470793
000d8313
00f12a23
00072d83
000217b7
88c78793
02f12a23
00000913
002a6a93
00200793
07800493
00000693
0cd103a3
fff00693
1ed30463
012de6b3
f7fafa13
1c069c63
24031263
18079e63
001afb93
1b010b13
1e0b90e3
0c714783
000b8a93
006bd463
00030a93
00012823
02012423
02012223
00012e23
ee0796e3
8edff06f
00044483
06800793
32f482e3
040a6a13
85dff06f
02b00793
00044483
0cf103a3
84dff06f
00044483
080a6a13
841ff06f
00044483
00140713
01749463
6850106f
fd048693
00070413
00000d93
82dae2e3
00044483
002d9793
01b787b3
00179793
00d78db3
fd048693
00140413
fedaf2e3
801ff06f
00044483
001a6a13
ff0ff06f
0c714783
00044483
fe079263
02000793
0cf103a3
fd8ff06f
000d8313
010a6a13
020a7793
080784e3
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
bffa7a93
00000793
eddff06f
000d8313
010a6a93
020af793
080780e3
01412783
00778b13
ff8b7b13
008b0793
00f12a23
000b2d83
004b2903
00100793
ea9ff06f
00044483
008a6a13
f60ff06f
000d8313
010a6a13
020a7793
7a078e63
01412783
00778b13
ff8b7b13
004b2783
000b2d83
008b0713
00e12a23
00078913
7c07c663
fff00793
000a0a93
02f30463
012de7b3
f7fa7a93
00079e63
02031263
000a8a13
00000313
00000b93
1b010b13
e69ff06f
2c091ce3
00900793
2db7e8e3
030d8d93
1bb107a3
000a8a13
00100b93
1af10b13
e45ff06f
000a0a93
00100693
fcd78ae3
00200693
06d78c63
1b010b13
01d91713
007df793
003ddd93
03078793
01b76db3
00395913
fefb0fa3
012de733
000b0613
fffb0b13
fc071ce3
001af693
06068a63
03000693
06d78663
ffe60613
1b010793
fedb0fa3
40c78bb3
000a8a13
00060b13
dd5ff06f
00100713
00e79463
3410106f
00200713
000a0a93
f8e798e3
03412683
1b010b13
00fdf793
00f687b3
0007c703
004ddd93
01c91793
01b7edb3
00495913
feeb0fa3
012de7b3
fffb0b13
fc079ce3
1b010793
41678bb3
000a8a13
d79ff06f
06500713
9e975ce3
0f012703
0a010593
0b010513
0ae12823
0f412703
04f12023
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
7ec0f0ef
04012783
40051463
0e812703
000216b7
8bc68693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
2ee6c6e3
0cc12703
02012683
6ad75063
03012703
02c12683
008c8c93
feecac23
0e812703
00d787b3
fedcae23
00170713
0ef12623
0ee12423
00700693
7ee6c663
02012703
fff70493
e8905463
01000693
0e812703
2a96dce3
01000913
00700b93
00c0006f
ff048493
2a9952e3
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
3a40b0ef
1c051463
0ec12783
0e812703
10c10c93
fb5ff06f
41598933
df205063
01000613
0e812703
09265463
04812023
01000e13
000c0413
00700d93
00090c13
00030913
00c0006f
ff0c0c13
058e5a63
00812683
01078793
00170713
00dca023
01cca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
00040593
000d0513
3240b0ef
20051ce3
01000e13
ff0c0c13
0ec12783
0e812703
10c10c93
fb8e4ae3
00090313
000c0913
00040c13
04012403
00812683
012787b3
00170713
00dca023
012ca223
0ef12623
0ee12423
00700693
008c8c93
d2e6d463
0e410613
000c0593
000d0513
04612023
2bc0b0ef
0e051063
0ec12783
04012303
10c10c93
d00ff06f
01000613
0e812703
07b65463
01000313
00700913
00c0006f
ff0d8d93
05b35a63
00812683
01078793
00170713
00dca023
006ca223
0ef12623
0ee12423
008c8c93
fce95ce3
0e410613
000c0593
000d0513
2540b0ef
06051c63
01000313
ff0d8d93
0ec12783
0e812703
10c10c93
fbb34ae3
00812683
01b787b3
00170713
00dca023
01bca223
0ef12623
0ee12423
00700693
008c8c93
c6e6d863
0e410613
000c0593
000d0513
2000b0ef
02051263
0ec12783
10c10c93
c50ff06f
0e410613
000c0593
000d0513
1e00b0ef
c8050a63
01012583
cc058063
000d0513
73c020ef
cb4ff06f
01000613
0e812703
00d64463
5e00106f
00020637
e2460d93
05212623
04812823
000d8913
000d0413
000a8d93
01000e13
00098a93
00700293
00048993
05f12023
000c0493
00068d13
000b0c13
00030b13
00c0006f
ff0d0d13
05ae5a63
01078793
00170713
012ca023
01cca223
0ef12623
0ee12423
008c8c93
fce2dee3
0e410613
00048593
00040513
13c0b0ef
7c051c63
01000e13
ff0d0d13
0ec12783
0e812703
10c10c93
00700293
fbae4ae3
000b0313
000d0693
000c0b13
00040d13
00048c13
04012f83
00098493
05012403
000a8993
000d8a93
00090d93
04c12903
00d787b3
00170713
00dca223
01bca023
0ef12623
0ee12423
00700693
008c8c93
aae6d663
0e410613
000c0593
000d0513
04612623
05f12023
0b00b0ef
ec051ae3
0ec12783
04c12303
04012f83
10c10c93
a7cff06f
0e410613
000c0593
000d0513
04612023
0840b0ef
ea0514e3
0ec12783
04012303
10c10c93
ac0ff06f
0cc12603
64c05e63
01c12703
02012683
00070493
38e6ce63
02905663
0e812703
009787b3
016ca023
00170713
009ca223
0ef12623
0ee12423
00700693
008c8c93
56e6c4e3
fff4c713
41f75713
00e4f4b3
01c12703
409704b3
44904663
01c12683
400a7713
00db04b3
0c0714e3
0cc12683
02012703
00e6c663
001a7713
54070ae3
03012703
02c12603
008c8c93
feecac23
0e812703
00c787b3
feccae23
00170713
0ef12623
0ee12423
00700613
00e65463
3b00106f
02012703
00eb0833
40d70633
40980933
01265463
00060913
03205863
0e812703
012787b3
009ca023
00170713
012ca223
0ef12623
0ee12423
00700693
008c8c93
00e6d463
3e80106f
fff94713
41f75713
00e97933
412604b3
9e905863
01000693
0e812703
6296d063
01000913
00700b93
00c0006f
ff048493
60995663
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
70d0a0ef
d20518e3
0ec12783
0e812703
10c10c93
fb5ff06f
001a7613
c4061663
00eca223
0ef12623
0e912423
00700713
ce975a63
0e410613
000c0593
000d0513
6cd0a0ef
ce0518e3
0ec12783
0e812483
10c10d93
cd0ff06f
cd205663
01000713
65275463
01000b93
00700b13
00c0006f
ff090913
632bda63
00812703
01078793
00148493
00eda023
017da223
0ef12623
0e912423
008d8d93
fc9b5ce3
0e410613
000c0593
000d0513
6650a0ef
c80514e3
0ec12783
0e812483
10c10d93
fb5ff06f
01412703
010a7793
00072d83
00470713
00e12a23
10079463
040a7793
0e078c63
010d9d93
410ddd93
41fdd913
00090793
8207dee3
01b037b3
41200933
40f90933
41b00db3
000a0a93
02d00693
00100793
e84ff06f
01412703
010a7793
00072d83
00470713
00e12a23
0a079263
040a7793
08078a63
010d9d93
010ddd93
00000913
f6cff06f
01412703
010af793
00072d83
00470713
00e12a23
06079063
040af793
04078663
010d9d93
010ddd93
00000913
00100793
e1cff06f
001a7713
00071463
81cff06f
959ff06f
000d8313
f74ff06f
00044483
00f12a23
ebdfe06f
03000793
1af107a3
1af10b13
e18ff06f
200af793
00078463
0ffdfd93
00000913
00100793
dd0ff06f
200a7793
300790e3
00000913
edcff06f
200a7793
2c0798e3
41fdd913
00090793
f44ff06f
03c12783
00044483
00079463
e61fe06f
0007c783
00079463
e55fe06f
400a6a13
e4dfe06f
00c12603
0006a783
00e12a23
41f65693
00c7a023
00d7a223
00040b13
fbdfe06f
01412703
00072783
00470713
00e12a23
0007a603
0047a683
0087a703
00c7a783
904ff06f
00068493
c69044e3
c8dff06f
000d8313
000a0a93
e5cff06f
000217b7
88c78793
000d8313
02f12a23
020a7793
12078863
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
001a7793
00078e63
012de7b3
00078a63
03000793
0cf10423
0c9104a3
002a6a13
bffa7a93
00200793
cccff06f
000217b7
8a078793
000d8313
02f12a23
fa1ff06f
000d8313
da8ff06f
00144483
020a6a13
00140413
d65fe06f
0e410613
000c0593
000d0513
40d0a0ef
a20518e3
0ec12783
10c10c93
ffcff06f
00144483
200a6a13
00140413
d35fe06f
00600793
000d8b93
13b7eee3
00021837
000b8a93
01212a23
8b480b13
d7dfe06f
01000693
0e812703
4296de63
01000b93
00700d93
00c0006f
ff048493
429bd463
00812683
01078793
00170713
00dca023
017ca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
000c0593
000d0513
3790a0ef
98051ee3
0ec12783
0e812703
10c10c93
fb5ff06f
01412703
010a7793
00072d83
00470713
00e12a23
06079663
040a7793
04078e63
010d9d93
010ddd93
00000913
ec5ff06f
0e410613
000c0593
000d0513
3250a0ef
940514e3
0ec12783
0e812483
10c10d93
884ff06f
0e410613
000c0593
000d0513
3010a0ef
920512e3
0ec12783
0e812483
10c10d93
88cff06f
200a7793
08079ae3
00000913
e6dff06f
1b010b13
00000793
00812823
00912e23
000b0413
03312223
000c0b13
000d8493
00090993
03c12d83
400afa13
0ff00b93
00030c13
00078913
0240006f
00a00613
00000693
00048513
00098593
36c0e0ef
52098c63
00050493
00058993
00a00613
00000693
00048513
00098593
10d0e0ef
03050513
fea40fa3
00190913
fff40413
fa0a0ee3
000dc683
fad91ae3
fb7908e3
4a099c63
00900793
4a97e863
000c0313
1b010793
000b0c13
00040b13
01c12483
02412983
01012403
03b12e23
03212023
41678bb3
000a8a13
ac4ff06f
0e812703
000216b7
8bc68693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
48e6cc63
18061c63
02012683
001a7713
00d76733
00071463
c55fe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
76e6ce63
02012683
00170713
0168a023
00f687b3
00d8a223
0ef12623
0ee12423
00700693
00888c93
00e6c463
bf9fe06f
fa9fe06f
00040d13
00048c13
f80ff06f
0e410613
000c0593
000d0513
1490a0ef
f6051663
0ec12783
10c10c93
cfcff06f
00812683
009787b3
009ca223
00dca023
00170713
0ef12623
0ee12423
00700693
00e6c463
b9dfe06f
f51fe06f
00040c13
f2cff06f
0f012783
0a010593
0b010513
0af12823
0f412783
0a012023
0a012223
0af12a23
0f812783
0a012423
0a012623
0af12c23
0fc12783
0af12e23
6490e0ef
4e0540e3
0c714783
04700713
38975c63
00021837
88080b13
00012823
02012423
02012223
00012e23
f7fa7a13
00300a93
00300b93
00000313
00078463
848ff06f
a49fe06f
01412783
00040b13
0007a783
00e12a23
00c12703
00e7a023
b41fe06f
00812703
012787b3
00148493
00eda023
e55fe06f
000b0513
f4cfe0ef
00050b93
fd9fe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
5ee6ce63
e80650e3
ff000693
40c004b3
52d656e3
01000913
00700b93
00c0006f
ff048493
50995ce3
00812683
01078793
00170713
00d8a023
0128a223
0ef12623
0ee12423
00888893
fcebdce3
0e410613
000c0593
000d0513
7bc0a0ef
de051063
0ec12783
0e812703
10c10893
fb5ff06f
0fc12783
5607c463
0c714783
04700713
3e975ae3
00021837
88880b13
eddff06f
00812683
009787b3
00170713
00dca023
009ca223
0ef12623
0ee12423
00700693
008c8c93
f4e6d863
0e410613
000c0593
000d0513
7500a0ef
d6051a63
0ec12783
10c10c93
f30ff06f
02012703
02412b83
00812e23
00eb0733
05412023
05312623
03512223
02812983
03612423
03c12403
04412a03
04812a83
00700d93
01000913
000c8693
00070b13
080b8663
08099663
fff40413
fffb8b93
0e812703
014787b3
0156a023
00170713
0146a223
0ef12623
0ee12423
00868693
0eedcc63
00044603
409b0cb3
01965463
00060c93
03905663
0e812603
019787b3
0096a023
00160613
0196a223
0ef12623
0ec12423
0ecdc263
00044603
00868693
fffcc513
41f55513
00acf733
40e60cb3
01904c63
00c484b3
f60b9ee3
12098ee3
fff98993
f7dff06f
0e812603
01994863
0580006f
ff0c8c93
05995863
00812703
01078793
00160613
00e6a023
0126a223
0ef12623
0ec12423
00868693
fccddce3
0e410613
000c0593
000d0513
6200a0ef
c4051263
ff0c8c93
0ec12783
0e812603
10c10693
fb994ce3
00812703
019787b3
00160613
00e6a023
0196a223
0ef12623
0ec12423
1acdc4e3
00044603
00868693
00c484b3
f65ff06f
0e410613
000c0593
000d0513
5c80a0ef
be051663
0ec12783
10c10693
ef1ff06f
0e410613
000c0593
000d0513
5a80a0ef
bc051663
00044603
0ec12783
10c10693
f09ff06f
04412783
04812583
00000913
40f40433
00078613
00040513
3e9070ef
001dc583
00a00613
00000693
00b03833
00048513
00098593
010d8db3
6390d0ef
ad1ff06f
00900793
ac97e4e3
b0dff06f
0e410613
000c0593
000d0513
5380a0ef
b4051e63
0cc12603
0ec12783
10c10c93
b4dff06f
00021837
87c80b13
c6dff06f
00030693
00200613
0b010a93
0d010793
0cc10713
0dc10813
000a8593
000d0513
04612823
04d12623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
0bb12e23
3dd030ef
02812703
04700793
01c12f03
02012e83
02412e03
04c12683
05012303
00050b13
04f70ae3
04600793
00d50933
10f716e3
00054703
03000793
38f702e3
0a010b93
0cc12783
00f90933
000b8593
000a8513
00612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
0a012023
0a012223
0a012423
0a012623
7c80e0ef
01c12303
00090693
02050263
0dc12683
0126fe63
03000713
00168793
0cf12e23
00e68023
0dc12683
ff26e8e3
416687b3
02f12023
0cc12703
04700793
00e12e23
02812703
70f70863
02812703
04600793
0af704e3
01c12783
02812603
04100693
fff78b93
0d712623
0ff4f793
00000713
00d61863
00f78793
0ff7f793
00100713
0cf10a23
02b00793
000bda63
01c12783
00100b93
40fb8bb3
02d00793
0cf10aa3
00900793
1377d4e3
0e310a13
000a0913
00a00593
000b8513
d49fd0ef
03050793
fef90fa3
000b8513
00a00593
cb1fd0ef
000b8a93
06300793
00090d93
00050b93
fff90913
fd57c6e3
03050693
0ff6f693
ffed8793
fed90fa3
2f47f6e3
0d610713
0080006f
0007c683
00d70023
00178793
00170713
ff4798e3
0e510793
0d610713
41b787b3
00f707b3
0d410713
40e787b3
02f12c23
02012703
03812683
00100793
00d70bb3
14e7dee3
02c12783
00fb8bb3
04012783
fffbca93
41fada93
bff7fa13
100a6a13
015bfab3
02012423
02012223
00012e23
05812783
5e078e63
02d00793
0cf103a3
00000313
001a8a93
c8cfe06f
0e410613
000c0593
000d0513
2b80a0ef
8c051e63
0ec12783
10c10c93
a80ff06f
00600b93
ec4ff06f
02012703
00eb0833
40d70633
40980933
b1265e63
00060913
b14ff06f
01412783
00e12a23
00c12703
0007a783
00040b13
00e79023
d40fe06f
018d9d93
418ddd93
41fdd913
00090793
c71fe06f
0ffdfd93
00000913
dd8ff06f
0ffdfd93
00000913
bddfe06f
02d00793
0cf103a3
a99ff06f
0e410613
000c0593
000d0513
2200a0ef
d08fe06f
0e410613
000c0593
000d0513
20c0a0ef
00050463
82cff06f
0cc12603
0ec12783
0e812703
10c10893
860650e3
9e1ff06f
05800793
03000713
0ce10423
002a6713
0cf104a3
04e12023
06300793
00012823
14c10b13
7c67c663
0fc12d83
fdf4f793
02f12423
04012c23
0f012e03
0f412e83
0f812f03
102a6a13
520dca63
06100793
00f48463
e78fe06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
578110ef
0cc10613
2c0070ef
00058613
00050593
000a8513
368110ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
7cc0e0ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
42c0e0ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000217b7
88c78793
02f12223
fff30913
06912023
07312423
07912823
07a12a23
07812c23
01c12483
00090c13
04812e23
07412223
06612623
000b0c93
07612e23
00068d13
000e0d93
000e8913
000f0993
0480006f
000b8593
000a8513
02c12023
01f12e23
0bf12c23
0ac12e23
0b612823
0b412a23
0a012023
0a012223
0a012423
0a012623
3840e0ef
fffc0c13
00090f93
00098613
0e050263
400307b7
00048613
000b8593
000a8513
08f12e23
0ba12023
0bb12223
0b212423
0b312623
08012823
08012a23
08012c23
6940e0ef
000a8513
76d100ef
00050593
00050413
000a8513
0b012a03
0b412983
0b812b03
0bc12903
060110ef
0b012683
04c12603
00048593
08d12023
0b412683
000b8513
09412823
08d12223
0b812683
09312a23
09612c23
08d12423
0bc12683
09212e23
08d12623
1f10f0ef
02412783
0a012b03
0a412a03
008786b3
0006c683
0a812f83
0ac12603
05912a23
00dc8023
05812823
fff00793
001c8c93
000b0d13
000a0d93
000f8913
00060993
eefc10e3
06c12303
000b0393
000a0293
3ffe0937
000b8593
000a8513
02612023
00812e23
06012483
05c12403
06412a03
0a712823
06712223
0a512a23
06512023
0bf12c23
05f12e23
0ac12e23
04c12623
0a012023
0a012223
0a012423
0b212623
3000e0ef
000c8d93
06812983
07012c83
07412d03
07812c03
07c12b03
02012303
44a04663
000b8593
000a8513
2080e0ef
02012303
00051863
01c12783
0017f913
42091663
05012783
03000693
00178713
00ed8733
0007c863
001d8d93
fedd8fa3
ffb71ce3
416d87b3
02f12023
a39ff06f
00130693
00200613
941ff06f
00030693
00300613
935ff06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
224110ef
0cc10613
76d060ef
00058613
00050593
000a8513
014110ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
4780e0ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
0d80e0ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000217b7
8a078793
02f12223
cadff06f
02812b03
02012703
02812e23
04012a03
00eb0733
01c12403
04c12983
02412a83
00068c93
00976463
d0dfe06f
00070493
d05fe06f
01c12703
ffd00793
00f74463
02e35463
ffe48493
fdf4f793
02f12423
8e5ff06f
0c714783
00000313
00078463
c94fe06f
e95fd06f
02012783
01c12703
1af74863
04012783
01c12703
0017f793
00070b93
00078663
02c12783
00f70bb3
04012783
4007f793
00078663
01c12783
2ef04863
fffbca93
41fada93
015bfab3
06700493
02012423
02012223
999ff06f
00012823
00078a13
800007b7
01b7cdb3
02d00793
04f12c23
ac1ff06f
04012783
00d50933
0017f793
0a079c63
0dc12683
81dff06f
0e410613
000c0593
000d0513
435090ef
00050463
a55fe06f
00044603
0ec12783
10c10693
00c484b3
da4ff06f
07800793
a2dff06f
0e410613
000c0593
000d0513
401090ef
00050463
a21fe06f
0cc12683
0ec12783
10c10c93
c31fe06f
02d00793
0cf103a3
b20ff06f
00020637
e2460d93
ae9fe06f
0c714783
01212a23
02012423
02012223
00012e23
00030a93
00030b93
00000313
00078463
b68fe06f
d69fd06f
00021837
88480b13
aecff06f
0a010b93
f0cff06f
0e410613
000c0593
000d0513
381090ef
00050463
9a1fe06f
0cc12483
02012703
0ec12783
10c10c93
40970633
bf1fe06f
04012783
01c12703
0017f793
0067e7b3
2ae05463
22079263
01c12b83
06600493
04012783
4007f793
18079a63
fffbca93
41fada93
015bfab3
ea5ff06f
000206b7
e2468d93
9f0fe06f
02012783
02c12703
06700493
00e78bb3
01c12783
fcf042e3
40fb8bb3
001b8b93
fffbca93
41fada93
015bfab3
e69ff06f
fff00793
00f12623
dd9fd06f
00812683
009787b3
00170713
00d8a023
0098a223
0ef12623
0ee12423
00700693
00888893
92e6d263
0e410613
000c0593
000d0513
2a5090ef
00050463
8c5fe06f
0ec12783
0e812703
10c10893
8fcff06f
0d610793
00071863
03000793
0cf10b23
0d710793
1b010713
030b8b93
40e78733
01778023
0dd70793
02f12c23
f3cff06f
05412783
000d8713
0cf12e23
02412783
fffdc683
00f7c603
02d61063
03000593
feb70fa3
0dc12703
fff70793
0cf12e23
fff74683
fed606e3
00168613
03900593
0ff67613
00b68663
fec70fa3
badff06f
02412783
00a7c603
fec70fa3
b9dff06f
00130593
000d0513
00612823
798040ef
01012303
00050b13
1a050663
00a12823
819ff06f
000a0a93
c2cfe06f
00030463
e81fd06f
00100313
e79fd06f
00600313
e71fd06f
04012783
0017f793
ea078463
e9cff06f
06700493
03c12603
0ff00713
00064783
14e78a63
01c12683
00000513
00000593
00d7de63
40f686b3
00164783
04078463
00158593
00160613
fee794e3
02c12e23
00d12e23
02b12223
02a12423
02812783
02412703
04412583
00e78533
a4cfd0ef
01750bb3
fffbca93
41fada93
015bfab3
e54ff06f
00064783
00150513
fbdff06f
02c12783
06600493
00f70bb3
006b8bb3
dd9ff06f
0a010b93
000b8593
000a8513
04612623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
04d12823
0bb12e23
0a012023
0a012223
0a012423
0a012623
4410d0ef
01c12f03
02012e83
02412e03
04c12303
c2050863
05012683
00100793
40d787b3
0cf12623
c20ff06f
00079a63
00100a93
06600493
00100b93
c15ff06f
02c12783
06600493
00178b93
006b8bb3
fffbca93
41fada93
015bfab3
bf5ff06f
00200793
02f12c23
d48ff06f
01412783
0007ad83
00478793
000dd463
fff00d93
00144483
00f12a23
00070413
98dfd06f
02012423
02012223
ee1ff06f
00cc5783
0407e793
00fc1623
b15fd06f
04007737
00050793
67472503
00060693
00058613
00078593
f98fd06f
00c5d783
0645ae03
00e5d303
01c5a883
0245a803
b8010113
ffd7f793
40000713
46812c23
00f11a23
00058413
07010793
00810593
46912a23
47212823
46112e23
00050913
07c12623
00611b23
03112223
03012623
00f12423
00f12c23
00e12823
00e12e23
02012023
f2cfd0ef
00050493
02055c63
01415783
0407f793
00078863
00c45783
0407e793
00f41623
47c12083
47812403
47012903
00048513
47412483
48010113
00008067
00810593
00090513
6a4000ef
fc0500e3
fff00493
fb9ff06f
fe010113
00812c23
00912a23
01212823
00112e23
01312623
00050913
00058493
00060413
00050663
03852783
14078a63
00c41703
01842683
00877793
00d42423
01071693
0106d693
08078463
01042783
08078063
00002637
00c6f6b3
0ff4f993
0ff4f493
0a068063
00042703
01442683
40f707b3
0ad7de63
00842683
00170613
00c42023
fff68693
00d42423
01370023
01442703
00178793
0cf70863
00c45783
0017f793
00078663
00a00793
0af48e63
01c12083
01812403
01012903
00c12983
00048513
01412483
02010113
00008067
00040593
00090513
0c8000ef
08051e63
00c41703
00002637
0ff4f993
01071693
0106d693
00c6f6b3
01042783
0ff4f493
f60694e3
06442683
00c76733
ffffe637
fff60613
00c6f6b3
00e41623
00042703
06d42223
01442683
40f707b3
f4d7c6e3
00040593
00090513
55c000ef
02051e63
00042703
00842683
00100793
00170613
fff68693
00c42023
00d42423
01370023
01442703
f2f71ce3
00040593
00090513
524000ef
f2050ee3
fff00493
f35ff06f
15d000ef
eadff06f
04007737
00050793
67472503
00058613
00078593
e65ff06f
040077b7
6747a783
ff010113
00812423
00912223
00112623
00050493
00058413
00078663
0387a703
08070463
00c41703
01071793
00877693
0107d793
08068863
01042683
0a068863
0017f613
02060863
01442603
00042423
00000513
40c00633
00c42c23
02068a63
00c12083
00812403
00412483
01010113
00008067
0027f613
00000593
00061463
01442583
00b42423
00000513
fc069ae3
0807f793
fc0786e3
04076713
00e41623
fff00513
fbdff06f
00078513
089000ef
00c41703
01071793
00877693
0107d793
f6069ce3
0107f693
08068263
0047f793
04079463
01042683
00876713
01071793
00e41623
0107d793
f4069ce3
2807f613
20000593
f4b606e3
00040593
00048513
7e1030ef
00c41703
01042683
01071793
0107d793
f2dff06f
03042583
00058e63
04040793
00f58863
00048513
1e5000ef
00c41703
02042823
01042683
fdb77713
00042223
00d42023
f91ff06f
00900793
00f4a023
04076713
00e41623
fff00513
f01ff06f
fd010113
000217b7
01412c23
a2c7aa03
03212023
02112623
148a2903
02812423
02912223
01312e23
01512a23
01612823
01712623
01812423
04090063
00050b13
00058b93
00100a93
fff00993
00492483
fff48413
02044263
00249493
009904b3
040b8463
1044a783
05778063
fff40413
ffc48493
ff3416e3
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
00492783
0044a683
fff78793
04878e63
0004a223
fa0688e3
18892783
008a9733
00492c03
00f777b3
02079263
000680e7
00492703
148a2783
01871463
f92784e3
f80788e3
00078913
f5dff06f
18c92783
0844a583
00f77733
00071c63
000b0513
000680e7
fcdff06f
00892223
fa9ff06f
00058513
000680e7
fb9ff06f
00c59783
fe010113
00812c23
01312623
00112e23
00912a23
01212823
0087f693
00058413
00050993
10069c63
00001737
80070713
0045a683
00e7e7b3
00f59623
18d05663
02842703
0c070c63
01079793
0107d793
000016b7
0009a483
00d7f6b3
0009a023
01c42583
16069863
00100693
00000613
00098513
000700e7
fff00793
18f50e63
00c45783
02842703
01c42583
0047f793
00078e63
00442683
03042783
40d50533
00078663
03c42783
40f50533
00050613
00000693
00098513
000700e7
fff00793
10f51e63
0009a703
00c41783
16070a63
01d00693
00d70663
01600693
0cd71463
01042683
fffff737
7ff70713
00e7f7b3
00f41623
00042223
00d42023
03042583
0099a023
00058c63
04040793
00f58663
00098513
770000ef
02042823
00000513
01c12083
01812403
01412483
01012903
00c12983
02010113
00008067
0105a903
fc090ee3
0005a483
01079713
01075713
00377713
0125a023
412484b3
00000793
00071463
0145a783
00f42423
00904863
fadff06f
00a90933
fa9052e3
02442783
01c42583
00048693
00090613
00098513
000780e7
40a484b3
fca04ee3
00c45783
fff00513
0407e793
01c12083
00f41623
01812403
01412483
01012903
00c12983
02010113
00008067
03c5a703
e6e04ae3
f4dff06f
05042503
eb5ff06f
00c45783
fffff737
7ff70713
00e7f7b3
01042683
01079793
4107d793
00c7d713
00f41623
00042223
00d42023
00177793
ee0788e3
04a42823
ee9ff06f
0009a783
e60782e3
01d00713
02e78863
01600713
02e78463
00c45783
0407e793
00f41623
ee5ff06f
fffff737
7ff70713
01042683
00e7f7b3
fa9ff06f
0099a023
00000513
ec5ff06f
fe010113
00812c23
00112e23
00050413
00050663
03852783
02078063
00c59783
02079663
01c12083
01812403
00000513
02010113
00008067
00b12623
40c000ef
00c12583
00c59783
fc078ee3
00040513
01812403
01c12083
02010113
d41ff06f
06050863
fe010113
040077b7
00812c23
00050413
6747a503
00112e23
00050663
03852783
02078a63
00c41783
00079c63
01c12083
01812403
00000513
02010113
00008067
00040593
01812403
01c12083
02010113
ce9ff06f
00a12623
38c000ef
00c41783
00c12503
fc0784e3
fd9ff06f
000217b7
a2c7a503
000075b7
7f458593
5b90006f
00000513
00008067
000125b7
e8858593
5a50006f
00000513
00008067
fe010113
000087b7
00112e23
00812c23
00912a23
01212823
01312623
01412423
01512223
01612023
00452403
8e078793
02f52e23
2ec50713
00300793
2ee52423
2ef52223
2e052023
00400793
00050913
00f42623
00800613
00000593
06042223
00042023
00042223
00042423
00042823
00042a23
00042c23
05c40513
a91fc0ef
0000eb37
00892483
0000eab7
0000ea37
0000e9b7
b90b0b13
bf4a8a93
c7ca0a13
ce498993
000107b7
03642023
03542223
03442423
03342623
00842e23
00978793
00f4a623
00800613
00000593
0604a223
0004a023
0004a223
0004a423
0004a823
0004aa23
0004ac23
05c48513
a21fc0ef
00c92403
000207b7
0364a023
0354a223
0344a423
0334a623
0094ae23
01278793
00f42623
06042223
00042023
00042223
00042423
00042823
00042a23
00042c23
05c40513
00800613
00000593
9d1fc0ef
01c12083
03642023
03542223
03442423
03342623
00842e23
01812403
00100793
02f92c23
01412483
01012903
00c12983
00812a03
00412a83
00012b03
02010113
00008067
ff010113
fff58793
00812423
00179413
00f40433
00241413
00f40433
00341413
01212023
00058913
07440593
00912223
00112623
3a9030ef
00050493
02050063
00c50513
0004a023
0124a223
00a4a423
06840613
00000593
931fc0ef
00c12083
00812403
00012903
00048513
00412483
01010113
00008067
fe010113
000217b7
01212823
a2c7a903
01312623
00112e23
03892783
00812c23
00912a23
01412423
00050993
0a078a63
2e090913
fff00493
00400a13
00492783
00892403
fff78793
0007d863
0840006f
06840413
06978e63
00c41703
fff78793
fe0718e3
ffff07b7
00178793
06042223
00042023
00042223
00042423
00f42623
00042823
00042a23
00042c23
00800613
00000593
05c40513
879fc0ef
02042823
02042a23
04042223
04042423
01c12083
00040513
01812403
01412483
01012903
00c12983
00812a03
02010113
00008067
00092403
00040c63
00040913
f61ff06f
00090513
d21ff0ef
f49ff06f
1ac00593
00098513
271030ef
00050413
02050663
00c50513
00042023
01442223
00a42423
1a000613
00000593
ff8fc0ef
00892023
00040913
f19ff06f
00092023
00c00793
00f9a023
f79ff06f
000217b7
a2c7a503
000125b7
e8858593
2550006f
03852783
00078463
00008067
cadff06f
00008067
00008067
00008067
00008067
040077b7
6747a503
000085b7
8d858593
17d0006f
040077b7
6747a503
000085b7
8ec58593
1690006f
ff010113
00812423
00000793
00000413
40f40433
00912223
00112623
40245493
02048063
ffc40413
00f40433
00042783
fff48493
ffc40413
000780e7
fe0498e3
00c12083
00812403
00412483
01010113
00008067
fe010113
01312623
040079b7
00812c23
00912a23
01212823
01412423
00112e23
00058a13
00050913
26498993
48c040ef
0089a703
000017b7
fef78413
00472483
41440433
ffc4f493
00940433
00c45413
fff40413
00c41413
00f44e63
00000593
00090513
461050ef
0089a783
009787b3
02f50863
00090513
444040ef
01c12083
01812403
01412483
01012903
00c12983
00812a03
00000513
02010113
00008067
408005b3
00090513
41d050ef
fff00793
04f50a63
040077b7
75078793
0007a703
0089a683
408484b3
0014e493
40870733
00090513
0096a223
00e7a023
3e0040ef
01c12083
01812403
01412483
01012903
00c12983
00812a03
00100513
02010113
00008067
00000593
00090513
3b9050ef
0089a703
00f00693
40e507b3
f4f6dce3
040076b7
6786a683
0017e793
00f72223
40d50533
040076b7
74a6a823
f39ff06f
12058a63
ff010113
00812423
00912223
00058413
00050493
00112623
35c040ef
ffc42803
ff840713
040075b7
ffe87793
00f70633
26458593
00462683
0085a503
ffc6f693
1ac50a63
00d62223
00187813
00d60533
0a081063
ff842303
00452803
04007537
40670733
00872883
26c50513
006787b3
00187813
14a88063
00c72303
0068a623
01132423
1e080463
0017e693
00d72223
00f62023
1ff00693
0af6e863
ff87f693
00868693
0045a503
00d586b3
0006a603
0057d813
00100793
010797b3
00a7e7b3
ff868513
00a72623
00c72423
00f5a223
00e6a023
00e62623
00812403
00c12083
00048513
00412483
01010113
28c0406f
00452503
00157513
02051e63
04007537
00d787b3
26c50513
00862683
0017e893
00f70833
16a68863
00c62603
00c6a623
00d62423
01172223
00f82023
f69ff06f
00008067
0017e693
fed42e23
00f62023
1ff00693
f4f6fce3
0097d693
00400613
0ed66c63
0067d693
03968813
03868613
00381813
01058833
00082683
ff880813
12d80863
0046a603
ffc67613
00c7f663
0086a683
fed818e3
00c6a803
01072623
00d72423
00812403
00c12083
00e82423
00048513
00412483
00e6a623
01010113
1c80406f
14081663
00c62583
00862603
00f686b3
00812403
00b62623
00c5a423
0016e793
00c12083
00f72223
00048513
00d70733
00412483
00d72023
01010113
1880406f
00187813
00d786b3
02081063
ff842503
40a70733
00c72783
00872603
00a686b3
00f62623
00c7a423
040077b7
0016e613
67c7a783
00c72223
00e5a423
eaf6e4e3
040077b7
78c7a583
00048513
c7dff0ef
e95ff06f
01400613
02d67463
05400613
06d66463
00c7d693
06f68813
06e68613
00381813
efdff06f
00d787b3
e99ff06f
05c68813
05b68613
00381813
ee5ff06f
00e5aa23
00e5a823
00a72623
00a72423
01172223
00f82023
e3dff06f
0045a503
40265613
00100793
00c797b3
00a7e7b3
00f5a223
ed5ff06f
15400613
00d66c63
00f7d693
07868813
07768613
00381813
e91ff06f
55400613
00d66c63
0127d693
07d68813
07c68613
00381813
e75ff06f
3f800813
07e00613
e69ff06f
0017e693
00d72223
00f62023
dcdff06f
00862783
32078063
00c5d683
fd010113
02812423
01412c23
01712623
02112623
02912223
03212023
01312e23
01512a23
01612823
01812423
01912223
01a12023
0086f793
00060b93
00050a13
00058413
08078663
0105a783
08078263
0026f793
000ba483
08078c63
02442783
01c42583
80000ab7
00000993
00000913
c00aca93
00098613
000a0513
04090263
00090693
012af463
000a8693
000780e7
26a05a63
008ba783
00a989b3
40a90933
40a787b3
00fba423
20078863
02442783
01c42583
00098613
000a0513
fc0912e3
0004a983
0044a903
00848493
fa9ff06f
00040593
000a0513
8f0ff0ef
3c051663
00c45683
000ba483
0026f793
f60798e3
0016f793
12079e63
00042783
00842703
80000ab7
ffeacb13
00000c13
00000993
fffaca93
00078513
00070c93
10098263
2006f613
24060e63
00070d13
2ee9ec63
4806f713
08070a63
01442603
01042583
00161713
00c70733
40b78933
01f75c93
00ec8cb3
00190793
401cdc93
013787b3
000c8613
00fcf663
00078c93
00078613
4006f693
2e068463
00060593
000a0513
39c030ef
00050d13
30050863
01042583
00090613
47d030ef
00c45783
b7f7f793
0807e793
00f41623
012d0533
412c87b3
01a42823
01942a23
00a42023
00098c93
00f42423
00098d13
000d0613
000c0593
569030ef
00842703
00042783
00098913
41970733
01a787b3
00e42423
00f42023
00000993
008ba783
012c0c33
412787b3
00fba423
0a078a63
00042783
00842703
00c45683
00078513
00070c93
f00992e3
0004ac03
0044a983
00848493
ee9ff06f
00000a93
00000513
00000c13
00000993
0e098063
0e050863
000a8793
00098b13
0137f463
00078b13
00042503
01042783
00842903
01442683
00a7f663
00d90933
0f694263
1adb4e63
02442783
01c42583
000c0613
000a0513
000780e7
00050913
06a05a63
412a8ab3
00100513
040a8c63
008ba783
012c0c33
412989b3
412787b3
00fba423
f80796e3
00000513
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00012d03
03010113
00008067
00040593
000a0513
bc0ff0ef
fa0500e3
00c41783
0407e793
00f41623
fff00513
fa9ff06f
00000513
00008067
0044a983
00048793
00848493
fe098ae3
0007ac03
00098613
00a00593
000c0513
209030ef
14050463
00150513
41850ab3
ef9ff06f
000c0593
00090613
3dd030ef
00042783
00040593
000a0513
012787b3
00f42023
b48ff0ef
f0050ee3
f89ff06f
01042683
04f6e863
01442903
0529e463
00098513
013b7463
000a8513
00090593
cf9fb0ef
00090593
ccdfb0ef
02442783
01c42583
00050693
000c0613
000a0513
000780e7
00050913
f2a05ee3
412989b3
e25ff06f
00070913
00e9f463
00098913
00078513
00090613
000c0593
34d030ef
00842703
00042783
41270733
012787b3
00e42423
00f42023
fc0712e3
00040593
000a0513
aa8ff0ef
ee0516e3
412989b3
dd5ff06f
00098c93
00098d13
d9dff06f
000b0613
000c0593
301030ef
00842703
00042783
000b0913
41670733
016787b3
00e42423
00f42023
e3dff06f
000a0513
6a9040ef
00050d13
d40510e3
01042583
000a0513
86dff0ef
00c41783
00c00713
00ea2023
f7f7f793
e81ff06f
00198793
00078a93
db9ff06f
00c00713
00c41783
00ea2023
e65ff06f
fff00513
e11ff06f
fe010113
01212823
01312623
01412423
01512223
01612023
00112e23
00812c23
00912a23
00058b13
2e050a93
00000a13
00100993
fff00913
004aa483
008aa403
fff48493
0204c663
00c45783
fff48493
00f9fc63
00e41783
00040513
01278663
000b00e7
00aa6a33
06840413
fd249ee3
000aaa83
fc0a92e3
01c12083
01812403
01412483
01012903
00c12983
00412a83
00012b03
000a0513
00812a03
02010113
00008067
fd010113
03212023
01312e23
01412c23
01512a23
01612823
01712623
02112623
02812423
02912223
00050a93
00058b93
2e050b13
00000a13
00100993
fff00913
004b2483
008b2403
fff48493
0204c863
00c45783
fff48493
00f9fe63
00e41783
00040593
000a8513
01278663
000b80e7
00aa6a33
06840413
fd249ce3
000b2b03
fc0b10e3
02c12083
02812403
02412483
02012903
01c12983
01412a83
01012b03
00c12b83
000a0513
01812a03
03010113
00008067
00450693
00000793
01a50513
ffff8837
01c0006f
00179793
00e69023
01079793
00268693
0107d793
02d50e63
0006d703
00177613
00060463
0017e793
00175713
0027f613
010765b3
fc0606e3
00179793
00b69023
01079793
00268693
0107d793
fcd516e3
00008067
01850693
00000713
00250513
01c0006f
00171713
00f69023
01071713
ffe68693
01075713
04d50463
0006d783
01079613
41065613
00179793
00065463
00176713
01079793
0107d793
00277613
0017e593
fc0600e3
00171713
00b69023
01071713
ffe68693
01075713
fcd510e3
00008067
fc010113
03312623
000109b7
02812c23
02912a23
03212823
03412423
03512223
02112e23
00050a13
00060493
00011d23
00011e23
01858913
01c10413
00810a93
fff98993
00095503
000a0593
ffe40413
ffe90913
02050a63
93dfb0ef
00245703
00045683
013577b3
00e787b3
01055513
0107d713
00d50533
00e50533
00a41023
00f41123
01055513
fea41f23
fb541ce3
00448613
01e10713
00045783
00240413
00260613
fef61f23
fee418e3
03c12083
03812403
03412483
03012903
02c12983
02812a03
02412a83
04010113
00008067
00055703
00255783
00070663
00008737
00e7e7b3
00f59923
00255703
000087b7
fff78793
02f70463
00650793
01058593
01850513
0007d703
00278793
ffe58593
00e59123
fea798e3
00008067
00650793
01a50513
0007d703
00278793
02071a63
fea79ae3
01258713
00058793
00278793
fe079f23
fef71ce3
0125d783
00008737
fff70713
00e7e7b3
00f59923
00008067
01058713
00058793
00278793
fe079f23
fef71ce3
ffffc7b7
00f59823
ffff87b7
fff7c793
00f59923
00008067
00455783
ff010113
00912223
00112623
00812423
01212023
00050493
0c079c63
00655703
00000413
01071793
4107d793
0a07c463
01a50693
0a000613
02071863
00648793
0080006f
0007d703
00278793
fee79e23
fed79ae3
00049c23
01040413
06c40c63
0064d703
fc070ce3
f0077793
04079063
01848513
00248593
00000793
00050713
00075683
ffe70713
00869613
00c7e7b3
00f71123
0086d793
feb714e3
0064d703
00840413
f0077793
fc0788e3
0a000913
0140006f
00140413
d49ff0ef
00894c63
0064d703
01071713
41075713
00048513
fe0752e3
00c12083
00040513
00812403
00412483
00012903
01010113
00008067
f007f713
00000413
04071063
f6f00913
0140006f
fff40413
c91ff0ef
fd2404e3
0044d783
00048513
fe0796e3
00c12083
00040513
00812403
00412483
00012903
01010113
00008067
00450693
01a50593
00000713
0080006f
0006d783
0087d613
00c76733
00879793
00e69023
01079713
00268693
01075713
fed590e3
0044d783
ff800413
f89ff06f
fe010113
00812c23
00912a23
00112e23
01212823
01312623
00058493
00050413
0a05c463
00f00793
00058613
00450513
01840693
00f00593
0297d463
00050793
0027d703
00278793
fee79f23
fef69ae3
00041c23
ff060613
fec5c2e3
00f4f493
00700793
0297d863
01840713
00240593
00000793
00075683
ffe70713
00869613
00c7e7b3
00f71123
0086d793
fee594e3
ff848493
00048a63
fff48493
00040513
be9ff0ef
fe049ae3
01c12083
01812403
01412483
01012903
00c12983
00000513
02010113
00008067
ff100793
40b00933
08f5de63
01850593
00000993
00450693
00f00613
01845703
00058793
00e9e9b3
ffe7d703
ffe78793
00e79123
fed79ae3
00041223
ff090913
fd264ee3
ff000913
ff100713
40990933
00000793
08e4ce63
00f90933
00700793
0527ca63
02090063
01845783
fff90913
00040513
0017f793
00f9e9b3
addff0ef
fe0914e3
01c12083
01812403
01412483
01012903
01303533
00c12983
02010113
00008067
ff900793
00000993
00450693
faf5dce3
01844783
01a40593
00f9e9b3
00000793
0006d703
00268693
00875613
00c7e7b3
00871713
fef69f23
01071793
0107d793
feb690e3
ff890913
f79ff06f
ff097793
40f007b3
00f90933
00700793
f727d2e3
fb1ff06f
01255783
00008637
fff60613
00f7d793
40f007b3
00f59023
01255683
01050793
00458713
00c6f6b3
00d59123
02c68663
00658713
00059223
ffe50513
0007d683
ffe78793
00270713
fed71f23
fef518e3
00059c23
00008067
01255603
00d67633
00d61e63
01250813
00050693
0006d603
00268693
00061e63
ff069ae3
01a58593
00270713
fe071f23
fee59ce3
00008067
00658713
00059223
ffc50513
0007d683
ffe78793
00270713
fed71f23
fea798e3
00008067
01255783
fb010113
04812423
fff7c793
04112623
01179713
00058413
00071e63
01250693
00050793
0007d703
00278793
08071c63
fed79ae3
01245783
fff7c793
01179713
06070063
00810593
f01ff0ef
02410593
00040513
ef5ff0ef
00815583
02415503
06b50c63
00a10793
02610713
02010613
0007d683
00278793
0a069863
00075683
00270713
0a069263
fef614e3
00000513
04c12083
04812403
05010113
00008067
00040793
0007d703
01240693
00278793
00071a63
f8d788e3
0007d703
00278793
fe070ae3
04c12083
04812403
ffe00513
05010113
00008067
00a15603
02615683
00153513
00a10713
02610793
00151513
fff50513
03c10593
00278793
00270713
00d61e63
f8b784e3
00075603
0007d683
00270713
00278793
fed606e3
f6c6eae3
40a00533
f6dff06f
00100513
f60582e3
fff00513
f5dff06f
fd010113
02812423
03212023
01312e23
01412c23
01512a23
01712623
00078913
00068b93
02112623
02912223
01612823
00050413
00058993
00060a13
00070a93
a85ff0ef
09000793
40ab8bb3
14a7d463
000087b7
ffe78793
2777d263
220a8c63
00492a83
00092683
01a90713
03490793
2ada8063
00270713
fe071f23
fee79ce3
03800793
32fa8263
1357d863
04000793
2afa8863
07100793
32fa9663
00008737
fff70713
000045b7
01400b13
00a00493
000087b7
00a00613
00860693
00169693
00e91a23
00992423
00b91b23
00f91c23
00c92623
00d90733
00f71523
01592023
01640b33
23705e63
000b5783
01495703
08f00693
00e7f633
0356cc63
00b00693
0296c863
00149713
00e40733
01840693
00275783
00078463
00166613
00071123
00270713
fee696e3
000b5783
01495703
fff74713
00e7f7b3
00fb1023
01695783
00c7f733
0c071463
13705263
00445783
22079663
000087b7
00041c23
ffe78793
1377cc63
01741123
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
03010113
00008067
160bd263
f7000793
12fbdc63
00240793
01a40413
00278793
fe079f23
fe879ce3
fb5ff06f
01800793
1afa8263
03500793
20fa9063
000017b7
7ff00713
40000593
00c00b13
00600493
80078793
00600613
ed5ff06f
01495703
000b5603
fff74793
00f677b3
00fb1023
01695783
00e67633
00c7f733
06070a63
02c79263
18099863
00c92783
01895703
00179793
00f407b3
0007d783
00e7f7b3
f0078ee3
03290513
01840613
01c90913
00000793
00055703
00065803
ffe60613
ffe50513
01070733
00f70733
01075793
00e61123
0017f793
fca91ee3
ef7042e3
09000793
00fa8663
00040513
e50ff0ef
00445783
0e079e63
00041c23
ec0bdee3
00041123
ed9ff06f
00041c23
ffff87b7
fff7c793
00f41123
00440793
01840413
00079023
00278793
fe879ce3
eb1ff06f
00240793
01a40413
00278793
fe079f23
fef41ce3
e99ff06f
000b8593
00040513
965ff0ef
00050463
00100993
d60a9ce3
00041c23
00041123
e75ff06f
e40a8ee3
00492a83
00092683
01a90713
03490793
d6da94e3
00892483
00149b13
01640b33
dd7046e3
09000793
ecfa82e3
01845783
00040513
0017f793
00f9e9b3
d28ff0ef
dadff06f
00010737
fff70713
000085b7
00e00b13
00700493
00100793
00600613
d5dff06f
0ff00713
08000593
00800b13
00400493
10000793
00400613
d41ff06f
00040513
ce0ff0ef
000087b7
001b8b93
00041c23
ffe78793
f177c2e3
ee0bcae3
dc9ff06f
e80a08e3
da5ff06f
0ff00713
08000593
00c00b13
00600493
10000793
00600613
cf9ff06f
00010737
fff70713
000085b7
01800b13
00c00493
00100793
00b00613
cd9ff06f
fd010113
03212023
01312e23
00058913
00255983
02112623
02812423
02912223
01412c23
00060493
01712623
01512a23
01612823
01812423
01912223
01a12023
00050b93
e9cff0ef
00295403
00050793
00090513
40f989b3
03448a13
e84ff0ef
40a40433
04e48713
000a0793
00278793
fe079f23
fee79ce3
09344863
004b8b13
00490a93
01ab8c13
00290d13
000a8713
000b0793
0007d603
00075683
00278793
00270713
0ad61a63
ff8796e3
018b8613
01890713
00000693
00075783
00065583
ffe70713
40d787b3
40b787b3
0107d693
00f71123
0016f693
ffe60613
fced1ee3
00100c93
000a0513
bfcff0ef
04c4d783
fff40413
00090513
00fce7b3
04f49623
be4ff0ef
f93454e3
00040693
02812403
02c12083
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00012d03
00048793
00090513
02412483
02012903
00000713
00000613
00000593
03010113
ac9ff06f
00000c93
f8c6e4e3
f4dff06f
fd010113
02812423
02112623
00058413
00410793
01e10713
00278793
fe079f23
fee79ce3
00e55603
000087b7
fff78793
00f65713
40e00733
00e11223
00f67633
06f60063
00e50793
00c11323
00a10713
ffe7d683
ffe78793
00270713
fed71f23
fef518e3
02061263
00011423
00040593
00410513
c4cff0ef
02c12083
02812403
03010113
00008067
00100793
fff00593
00410513
00f11423
e60ff0ef
fd1ff06f
00050793
00e50693
0007d703
00278793
06071c63
fef69ae3
01440713
00040793
00278793
fe079f23
fee79ce3
01240713
00040793
00278793
fe079f23
fef71ce3
01245783
000086b7
fff68693
00d7e7b3
01079793
0107d793
00f41923
00e51683
f606dce3
00040693
0006d603
00268693
f60614e3
fed71ae3
ffff8737
00e7c7b3
00f41923
f55ff06f
01040713
00040793
00278793
fe079f23
fee79ce3
ffffc7b7
00f41823
ffff87b7
fff7c793
00f41923
f29ff06f
01255783
f5010113
0a812423
fff7c793
0a912223
0b212023
09312e23
0a112623
09412c23
09512a23
09612823
09712623
09812423
09912223
09a12023
07b12e23
01179713
00050493
00058993
00060413
00068913
00071e63
01250693
00050793
0007d703
00278793
2e071a63
fed79ae3
0129d783
fff7c793
01179713
00071e63
01298693
00098793
0007d703
00278793
2e071463
fed79ae3
00020a37
e44a0593
00048513
f84ff0ef
2e050663
0124d603
0129d703
000087b7
fff78793
00f67533
00f775b3
0af51663
01248813
00048793
0007d683
00278793
08069863
ff079ae3
000087b7
fff78793
2cf59263
01298693
00098793
0007d583
00278793
48059663
fed79ae3
01040713
00040793
00278793
fe079f23
fee79ce3
ffffc7b7
00f41823
ffff87b7
fff7c793
00f41923
0ac12083
0a812403
0a412483
0a012903
09c12983
09812a03
09412a83
09012b03
08c12b83
08812c03
08412c83
08012d03
07c12d83
0b010113
00008067
000087b7
fff78793
24f58863
00048513
01c10593
df8ff0ef
03810593
00098513
decff0ef
03a15a83
01e15483
2a0a8e63
01512623
00048713
00912423
02010793
03410693
02071263
38d78c63
0007d703
00278793
fe070ae3
01c10513
a64ff0ef
40a487b3
00f12423
03812703
03890a93
000a8793
02e92a23
04e90493
00278793
fe079f23
fef49ce3
03810513
fd1fe0ef
02215b03
000109b7
05010c13
010b1a13
416a0a33
03a10c93
fff98993
06e10d13
05610d93
03c15503
03e15783
00098b93
01051513
00f50533
00aa6a63
000b0593
a25fa0ef
01051b93
010bdb93
05410613
01c10593
000b8513
84cff0ef
03c10713
05810793
0007d603
00075683
00278793
00270713
20d61a63
ffa796e3
00000793
06c10693
000c0613
00065703
0006d583
ffe60613
40f70733
40b70733
01075793
00e61123
0017f793
ffe68693
fd961ee3
017a9023
03c10793
0027d703
00278793
fee79f23
ff879ae3
04011823
002a8a93
f5549ae3
00000713
03c10793
05210613
0007d683
00278793
00d76733
fec79ae3
00e035b3
03810793
03490713
00075683
00278793
00270713
fed79f23
fef618e3
00c12783
00812703
000046b7
fff68693
40e78ab3
03810513
00090793
04000713
00da86b3
00000613
e34ff0ef
03815703
01c15783
00040593
03810513
40e787b3
00f037b3
40f007b3
02f11c23
818ff0ef
dd5ff06f
01448713
0004d783
00248493
00240413
fef41f23
fee498e3
db9ff06f
01440713
0009d783
00240413
00298993
fef41f23
fee418e3
d9dff06f
e44a0593
00098513
c8cff0ef
d00516e3
d61ff06f
dc0806e3
01440793
00240413
fe041f23
fef41ce3
d71ff06f
00000813
01298693
00098793
0007d583
00278793
fc059ae3
fed79ae3
000087b7
fff78793
04f50a63
00f65613
0009d783
00298993
18079263
fed99ae3
00f75793
00c7c7b3
00f79793
00f41923
01240713
00040793
00278793
fe079f23
fee79ce3
01245783
00008737
fff70713
00e7e7b3
00f41923
cf9ff06f
01248593
0004d783
00248493
12079e63
feb49ae3
f9dff06f
03c10793
05010c13
0cfc0e63
0007d703
00278793
fe070ae3
03810513
fbdfe0ef
40a007b3
01e15703
00f12623
d25ff06f
dec6fae3
fffb8793
01079513
01055513
00000693
03410613
06c10713
00075783
00065583
ffe70713
40d787b3
40b787b3
0107d693
00f71123
0016f693
ffe60613
fdb71ee3
03c10713
05810793
0007d603
00075683
00278793
00270713
00d61863
ffa796e3
00050b93
d8dff06f
fec6fce3
ffeb8893
01089b93
010bdb93
00000693
03410613
06c10713
00075783
00065583
ffe70713
40d787b3
40b787b3
0107d693
00f71123
0016f693
ffe60613
fdb71ee3
d45ff06f
01440793
00240413
fe041f23
fef41ce3
be9ff06f
01c15683
03815603
01240713
00040793
40c686b3
00d036b3
00f69693
00d41923
00278793
fe079f23
fef71ce3
eadff06f
00000793
e85ff06f
00000613
e69ff06f
00100813
e3dff06f
f7010113
08912223
00050493
01255503
00008737
fff70713
08812423
09212023
07412c23
08112623
07312e23
07512a23
07612823
07712623
07812423
07912223
00e57833
00058913
00060413
00068a13
00e81e63
01248993
00048713
00075603
00270713
1e061463
ff371ae3
01295603
000087b7
fff78793
00f675b3
08f58863
1ef81463
01248993
00048793
0007d703
00278793
26071663
fef99ae3
000205b7
e4458593
00090513
9f0ff0ef
22050463
01295603
000087b7
fff78793
00f675b3
24f58663
0124d503
00f57733
18f71e63
00048793
0007d703
00278793
3c071063
fef99ae3
0004d783
00248493
36079c63
ff349ae3
00f55713
000087b7
fff78793
0cf59063
01290693
0a80006f
01290693
00090713
00075783
00270713
18079e63
fee69ae3
000087b7
fff78793
f4f80ce3
00090793
0007d703
00278793
0e071863
fef69ae3
000205b7
e4458593
00048513
948ff0ef
18050063
0124d503
01295603
000087b7
fff78793
00f57833
00f675b3
0cf80a63
000087b7
fff78793
0ef59663
01290693
00090793
0007d703
00278793
0c071c63
fed79ae3
000087b7
fff78793
00f55713
00080593
01248993
f2f80ce3
00095783
00290913
2a079a63
fed91ae3
00f65793
00e7c7b3
00f79793
00f41923
01240713
00040793
00278793
fe079f23
fee79ce3
01245783
00008737
fff70713
00e7e7b3
00f41923
08c12083
08812403
08412483
08012903
07c12983
07812a03
07412a83
07012b03
06c12b83
06812c03
06412c83
09010113
00008067
0124d503
000087b7
fff78793
00f575b3
00058813
f4f592e3
01248993
e89ff06f
01440713
0004d783
00240413
00248493
fef41f23
fee418e3
f95ff06f
00048513
00c10593
f75fe0ef
02810593
00090513
f69fe0ef
00e15483
02a15983
08049663
01010793
02410693
1ef68063
0007d703
00278793
fe070ae3
00c10513
bf1fe0ef
02a15703
40a004b3
0640006f
01490713
00095783
00290913
00240413
fef41f23
fee918e3
f29ff06f
01040713
00040793
00278793
fe079f23
fee79ce3
ffffc7b7
00f41823
ffff87b7
fff7c793
00f41923
efdff06f
000087b7
fff78793
dcf594e3
01290693
e21ff06f
00098713
00098913
02c10793
04010693
02071263
16d78063
0007d703
00278793
fe070ae3
02810513
b5dfe0ef
02a15703
40a98933
02815783
038a0993
02ea1b23
02fa1a23
04ea0713
00098793
00079023
00278793
fee79ce3
04ca0c13
00000b93
02410a93
01010c93
04610b13
000ad503
ffea8a93
08051c63
04ca5783
000c0713
00fbebb3
ffe75603
ffe70713
00c71123
fee99ae3
020a1c23
fd9a9ae3
034a0713
02810793
04210613
00075683
00278793
00270713
fed79f23
fec798e3
ffffc6b7
012484b3
00268693
000b8593
02810513
000a0793
04000713
00d486b3
00000613
fe1fe0ef
02815703
00c15783
00040593
02810513
40e787b3
00f037b3
40f007b3
02f11423
9c5fe0ef
dddff06f
04410613
02810593
8e5fe0ef
000c0513
00000593
05c10613
00055783
00065703
ffe50513
ffe60613
00f70733
00b70733
01075593
00e51123
0015f593
fd661ee3
f2dff06f
00000713
c91ff06f
00000793
d55ff06f
01440793
00240413
fe041f23
fef41ce3
d75ff06f
01440793
00240413
fe041f23
fef41ce3
d61ff06f
00008837
fff80813
cd1ff06f
00c5a883
e1010113
0005ae83
0045ae03
0085a303
03112e23
04052583
fff00893
1e812423
17112023
00078413
09000893
09000793
1d412c23
1e112623
1e912223
1f212023
1d312e23
1d512a23
1d612823
1d712623
1d812423
1d912223
1da12023
1bb12e23
03d12823
03c12a23
02612c23
17112223
00c12023
00d12423
00e12823
01012a23
00f12623
00050a13
02058463
04452703
00100793
00e797b3
00f5a423
00e5a223
1e8020ef
16412783
040a2023
00f12623
06010913
00090593
03010513
bb4ff0ef
07215783
00008737
fff70713
00e7f5b3
00e59e63
00090713
07210613
00075683
00270713
3c0694e3
fec71ae3
00f7d793
00012703
00f42023
00300793
08f70ae3
01400793
00f12223
3a0716e3
000087b7
fff78793
00f59e63
00090793
07210693
0007d703
00278793
0e0712e3
fed79ae3
09000793
16f12223
07c10713
00090793
07410613
0007d683
00278793
00270713
fed71f23
fec798e3
08e15603
00012c23
01061793
4107d793
5607c863
00020bb7
e44b8d93
014d8c13
00000693
09810793
000c0713
0ac10d13
0080006f
00075683
00278793
fed79f23
00270713
ffa798e3
14060463
000087b7
fff78793
4af60ee3
08c11783
5207dce3
07c10593
000c0513
c2dfe0ef
12050e63
060542e3
08e15783
5c0796e3
08c11783
00000493
16010993
0207c463
118d8413
07c10613
00098693
00060593
00040513
95dff0ef
08c11783
fff48493
fe07d2e3
0d010413
0e810b13
00040713
07c10793
09010613
0007d683
00278793
00270713
fed71f23
fec798e3
00000693
09810793
000c0713
0080006f
00075683
00278793
fed79f23
00270713
ffa798e3
028d8d13
12cd8c93
fffffab7
21cd8d93
00c0006f
014c8c93
014d0d13
00040593
000c0513
b75fe0ef
04a05863
00040593
000c8513
b65fe0ef
02054863
00098693
00040613
00040593
000d0513
8b5ff0ef
09810613
00098693
00060593
000d0513
8a1ff0ef
015484b3
01fad793
015787b3
4017da93
fbbc90e3
09810613
00098693
000c0593
00060513
ae8ff0ef
12410a93
0300006f
07c10793
08e10693
0007d703
ec0712e3
00278793
fed79ae3
00000493
12410a93
16010993
0d010413
0e810b13
00040593
09810513
a1dfe0ef
09810713
00040793
0007d683
00278793
00270713
fed71f23
ff6798e3
00040593
07c10513
0a011823
9f1fe0ef
07c10793
00045703
00240413
00278793
fee79f23
ff6418e3
09810513
00098613
07c10593
08011a23
f99fe0ef
1ac15503
16051a63
09410c13
07e10c93
0b610413
e44b8593
07c10513
a59fe0ef
14050c63
00000713
000c0693
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fd9690e3
0b410713
07c10793
0007d683
00278793
00270713
fed71f23
ff8798e3
0c011623
00000713
0cc10693
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fc8690e3
00000713
0cc10693
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fc8690e3
00000613
000c0693
0cc10713
0006d583
00075783
ffe68693
ffe70713
00b787b3
00c787b3
0107d613
00f69123
00167613
fc871ee3
09810513
00098613
07c10593
e2dfe0ef
1ac15503
fff48493
ea0500e3
01812783
00012683
00300713
00f037b3
40f007b3
00d7f793
02078793
12f10223
00412783
00e69463
009787b3
02a00713
00f12c23
00f75463
00e12c23
00a00713
4ae50463
03050513
02e00713
12a102a3
12e10323
1c07c4e3
12710b13
00000413
00912e23
000b0493
00040b13
01812403
0b410c93
09410d13
07e10d93
0b610c13
00000693
000d0613
00065783
01079593
4105d593
0005d463
0016e693
00179793
01079793
0026f593
0107d793
00058463
0017e793
00169693
00f61023
01069693
ffe60613
0106d693
fdb610e3
000c8693
07c10793
0007d603
00278793
00268693
fec69f23
ffa798e3
0c011623
00000693
0cc10613
00065783
01079593
4105d593
0005d463
0016e693
00179793
01079793
0026f593
0107d793
00058463
0017e793
00169693
00f61023
01069693
ffe60613
0106d693
fd8610e3
00000693
0cc10613
00065783
01079593
4105d593
0005d463
0016e693
00179793
01079793
0026f593
0107d793
00058463
0017e793
00169693
00f61023
01069693
ffe60613
0106d693
fd8610e3
00000593
000d0613
0cc10693
00065503
0006d783
ffe60613
ffe68693
00a787b3
00b787b3
0107d593
00f61123
0015f593
fd869ee3
00098613
07c10593
09810513
c59fe0ef
1ac15603
00148793
001b0b13
03060693
fed78fa3
03644463
00078493
e9dff06f
01161613
000107b7
01165613
fff78793
08c11723
00f12c23
a7dff06f
00048b13
01c12483
00400713
04c75a63
00500713
00e60ae3
ffe7c703
01812683
ffe78613
07f77713
0206c663
02e00793
03800593
03000513
76f70663
78e5d263
fff64703
00a60023
fff60613
07f77713
fe9ff06f
03100713
fee78f23
00148493
000215b7
00048613
8dc58593
000b0513
3f8030ef
07215783
00c12703
16912823
fff7c793
16e12223
01179713
18070863
01012683
12414703
00148793
00f6a023
000a8793
02070a63
02e00693
20d70663
0017c703
00178793
fe071ae3
04500693
00fae663
0140006f
01578863
fff7c703
fff78793
fed71ae3
00078023
000a8793
02000693
02d00613
0007c703
00d70463
00c71663
00178793
ff1ff06f
000a8413
00c0006f
0007c703
00068413
00e40023
00140693
00178793
fe0716e3
00012703
00200793
fff44683
12f70063
00412783
00078713
0097d463
00048713
03000793
02f69663
415407b3
02f75263
03000693
00c0006f
415407b3
00f75a63
ffe44783
fe040fa3
fff40413
fed786e3
00012703
00300793
0ef70663
00812783
040a2223
00978613
01700793
10c7f663
00100713
00400793
00179793
01478693
00070593
00170713
fed678e3
04ba2223
000a0513
13d010ef
00050493
080502e3
04aa2023
000a8593
5f8030ef
01412703
00070863
415407b3
00f487b3
00f72023
1ec12083
1e812403
1e012903
1dc12983
1d812a03
1d412a83
1d012b03
1cc12b83
1c812c03
1c412c83
1c012d03
1bc12d83
00048513
1e412483
1f010113
00008067
00090793
07210693
0007d703
00278793
5a071063
fed79ae3
01012703
000027b7
70f78793
00f72023
e99ff06f
03000793
f2f696e3
415407b3
00100713
eef74ae3
f1dff06f
00412783
009784b3
4e04c063
01012783
00812703
0007a783
00f707b3
00f12423
00812783
040a2223
00378613
01700793
eec7eee3
00000593
f15ff06f
00812783
00078713
00f12223
02a00793
f6e7d663
00f12223
f64ff06f
0007c703
e00700e3
0017c703
00178793
fee78fa3
de0708e3
0017c703
00178793
fee78fa3
fe0712e3
dddff06f
03100713
12e102a3
02e00713
12e10323
00148493
2af05a63
03000793
12f103a3
01812783
12810b13
fff78793
00f12c23
b45ff06f
12410a93
000215b7
94858593
000a8513
000024b7
13c030ef
70f48493
d41ff06f
0b410c93
000c8713
07c10793
09010613
0007d683
00278793
00270713
fed71f23
fec798e3
000047b7
08e78793
0cf11323
000087b7
fff78793
00f12e23
ffffc7b7
12410a93
0d010413
01000713
0c8d8313
00278793
03412423
03512223
00000493
00040a93
16010993
0aa10b13
02f12023
00030a13
00070413
00098693
09810613
000c8593
000a0513
b11fe0ef
04c10713
09810793
0007d683
00278793
00270713
fed71f23
ffa798e3
01c12783
05e15583
00f5f533
02012783
00f50533
36a05463
09000613
40a60633
000a8713
04c10793
0007d683
00278793
00270713
fed71f23
ff2798e3
06c05663
00f00793
000a8713
02c7de63
08000693
40a686b3
0046d693
00168713
00171713
00ea8733
000a8793
00278793
fe079f23
fef71ce3
08000613
40a60633
00469693
40d60633
00161793
00fd87b3
00075683
2307d783
00f6f7b3
00f71023
01059593
4105d593
1405c463
09810793
000a8713
0007d603
00075683
02d61863
00278793
00270713
fefb16e3
000c8713
09810793
0007d683
00278793
00270713
fed71f23
ffa798e3
008484b3
014a0a13
12cd8793
00145413
ecfa1ee3
0c615783
08e15703
000a8413
02812a03
00e787b3
ffffc737
f7270713
02412a83
00e787b3
0cf11323
07c10713
000c8793
0c810613
0007d683
00278793
00270713
fed71f23
fec798e3
00000713
09810793
0080006f
000c5703
00278793
fee79f23
002c0c13
ffa798e3
028d8b13
00001c37
118d8d93
0100006f
001c5c13
25bb0463
014b0b13
000c8593
000d8513
994fe0ef
22a04a63
000c8593
000b0513
984fe0ef
fca04ce3
00098693
000c8613
000c8593
000b0513
945fe0ef
09810613
00098693
00060593
000b0513
ec1fe0ef
018484b3
fa9ff06f
12710b13
aa0798e3
8a5ff06f
00000793
c40ff06f
00812783
fff78793
cd9ff06f
04c10793
000a8713
0140006f
00278793
05e10693
00270713
ead782e3
0007d603
00075683
fed604e3
0e215783
01c12703
00e7f7b3
3ce78063
0ec10593
000c0513
838fe0ef
10810593
000a8513
82cfe0ef
0ec15703
10a15603
0ee15883
fff74713
01071713
01075713
0ee11623
40c885b3
00060693
06b05e63
02412583
10810693
12010793
0006d503
00268693
00258593
fea59f23
fef698e3
12011e23
10810693
0ec10593
0080006f
0005d703
00268693
fee69f23
00258593
fef698e3
02412783
12011023
0ec10713
13c10513
0007d683
00278793
00270713
fed71f23
fea798e3
10a15683
411605b3
10011223
00068613
32058c63
02d12623
f6f00793
06f5c863
0ec10513
da5fd0ef
02c12683
00050593
12010793
10410713
0ec15503
10815603
3ac50863
00000613
10a10893
00060513
0007d603
00075803
ffe78793
40a60633
41060633
01065513
00c79123
00157513
ffe70713
fd179ee3
00100613
00098793
04000713
10810513
900fe0ef
000a8593
10810513
afdfd0ef
d45ff06f
01012783
12010223
000a8413
0007a023
b29ff06f
000a8793
0e410713
00278793
fe079f23
fee79ce3
d0dff06f
01812783
12410a93
10078263
000215b7
8c058593
000a8513
000024b7
4d9020ef
70f48493
8ddff06f
0e810b13
c80ff06f
fff64783
03800713
0ef77863
03100793
00148493
fef60fa3
8a5ff06f
00170713
00e60023
899ff06f
07210713
0080006f
8ae90ee3
00095783
00290913
fe078ae3
01012703
000027b7
70f78793
00f72023
8e9ff06f
12410a93
000215b7
8d858593
000a8513
000024b7
45d020ef
70f48493
861ff06f
1ac15603
12610b13
12710793
fe4ff06f
09810593
07c10513
00f12e23
a09fd0ef
e44b8593
09810513
eb9fd0ef
01c12783
fc051863
01812703
800748e3
ffe7c703
fd270613
00163613
fff64613
00cb0633
00064603
00167613
fe060863
ffe78613
07f77713
fb0ff06f
000215b7
8cc58593
000a8513
000024b7
3d9020ef
70f48493
fdcff06f
00178793
fef60fa3
fbcff06f
0d010413
00040593
07c10513
00004cb7
d8dfd0ef
00000493
0e810b13
0cc10993
0d210a93
ffec8c93
0e815783
0077f793
0c079a63
0b410713
00040793
0007d683
00278793
00270713
fed71f23
ff6798e3
0b410513
0c011623
f94fd0ef
0b410513
f8cfd0ef
00000613
00098693
000b0713
0006d583
00075783
ffe68693
ffe70713
00b787b3
00c787b3
0107d613
00f69123
00167613
fd571ee3
0b615783
0b815703
00378793
0af11b23
02070063
0b410513
f3cfd0ef
0b615783
0b815703
00178793
0af11b23
fe0714e3
0cc15783
02079c63
0b615783
02fce863
00040713
0b410793
0007d683
00278793
00270713
fed71f23
ff3798e3
0e011423
fff48493
fd500793
f2f494e3
07c10593
00040513
889fd0ef
16010993
960ff06f
000a8793
0007d703
00278793
aa071ee3
0e210713
fee798e3
000a8793
0007d703
00278793
c20710e3
0e210713
fee798e3
a99ff06f
10c10713
0f010793
0007d883
00075503
00278793
00270713
04a89863
10610513
fea794e3
0ec15703
10815783
04f70663
000a8793
0e410713
00278793
fe079f23
fee79ce3
a51ff06f
000216b7
000015b7
00021537
8e068693
00000613
b6e58593
8f450513
30d060ef
07156c63
12010793
10410713
c7dff06f
00068713
00069663
10e11783
0c07d663
10a10713
12010793
00075583
10059663
00270713
fee79ae3
10c11523
ca1ff06f
00000613
0ee10893
0007d803
00075503
ffe78793
ffe70713
01050533
00c50633
01065513
00c79123
00157613
fd171ee3
00000613
c59ff06f
02412603
10810713
12010793
00075503
00270713
00260613
fea61f23
fef718e3
12011e23
10810513
0ec10613
10410713
00065803
00260613
00250513
ff051f23
fee618e3
02412603
12011023
0ec10893
13c10513
00065803
00260613
00288893
ff089f23
fea618e3
10011223
ba5ff06f
12010693
10a10893
0006d783
01079613
41065613
00065463
00176713
00179793
01079793
00277613
0107d793
00060463
0017e793
00171713
00f69023
01071713
ffe68693
01075713
fd1690e3
ba9ff06f
00168613
10c11523
b9dff06f
00852703
00c52783
00052603
00452683
fc010113
00010513
01410593
00e12423
00f12623
02112e23
00c12023
00d12223
9acfe0ef
02615783
00000513
fff7c793
01179713
02071063
01410793
02610693
0007d703
00278793
00071c63
fed79ae3
00200513
03c12083
04010113
00008067
00100513
ff1ff06f
0f050513
00008067
04007537
1e850513
00008067
04007537
1e850513
00008067
ff010113
00112623
00812423
00912223
02060c63
000215b7
95458593
00060513
00060413
1e5020ef
000214b7
02051263
95048513
00c12083
00812403
00412483
01010113
00008067
000214b7
fe5ff06f
95048593
00040513
1b1020ef
fc050ae3
000205b7
70c58593
00040513
19d020ef
fc0500e3
00000513
fbdff06f
040077b7
2207c503
00008067
ff010113
00112623
00812423
00912223
02058c63
00058413
000215b7
95458593
00040513
15d020ef
000214b7
02051263
95048513
00c12083
00812403
00412483
01010113
00008067
000214b7
fe5ff06f
95048593
00040513
129020ef
fc050ae3
000205b7
70c58593
00040513
115020ef
fc0500e3
00000513
fbdff06f
00c5d783
f8010113
06812c23
06112e23
06912a23
07212823
07312623
07412423
0027f713
00058413
02070c63
04358793
00f5a023
00f5a823
00100793
00f5aa23
07c12083
07812403
07412483
07012903
06c12983
06812a03
08010113
00008067
00e59583
00050493
0805cc63
00810613
5b1060ef
08054463
00c12783
0000f937
000019b7
00f97933
ffffe7b7
00f90933
00193913
40000a13
80098993
000a0593
00048513
1c8000ef
00c41783
06050e63
00008737
8e070713
02e4ae23
0807e793
00f41623
00a42023
00a42823
01442a23
08091863
0137e7b3
07c12083
00f41623
07812403
07412483
07012903
06c12983
06812a03
08010113
00008067
00c45783
0807f793
00000913
04078663
04000a13
000a0593
00048513
154000ef
00c41783
00000993
f80516e3
2007f713
f0071ae3
ffc7f793
0027e793
04340713
00f41623
00100793
00e42023
00e42823
00f42a23
ef1ff06f
40000a13
00000993
f41ff06f
00e41583
00048513
521060ef
00051663
00c41783
f61ff06f
00c45783
ffc7f793
0017e793
01079793
4107d793
f49ff06f
f9010113
06812423
00058413
00e59583
06912223
07212023
06112623
00060493
00068913
0405ca63
00810613
465060ef
04054463
00c12703
0000f7b7
06c12083
00e7f7b3
ffffe737
00e787b3
06812403
0017b793
00f92023
40000713
00e4a023
00001537
06412483
06012903
80050513
07010113
00008067
00c45783
0807f793
02078863
06c12083
06812403
00000793
00f92023
04000713
00e4a023
06012903
06412483
00000513
07010113
00008067
06c12083
06812403
00000793
00f92023
40000713
00e4a023
06012903
06412483
00000513
07010113
00008067
fd010113
01312e23
02112623
02812423
02912223
03212023
01412c23
01512a23
01612823
01712623
01812423
01912223
00b58793
01600713
00050993
06f76663
01000793
1eb7e663
2f5000ef
01000493
01800793
00200613
04007937
26490913
00f907b3
0047a403
ff878713
20e40a63
00442783
00c42683
00842603
ffc7f793
00f407b3
0047a703
00d62623
00c6a423
00176713
00098513
00e7a223
2a5000ef
00840513
1980006f
ff87f493
1807c263
18b4e063
289000ef
1f700793
4697f663
0094d793
1a078663
00400713
3cf76c63
0064d793
03978613
03878513
00361693
04007937
26490913
00d906b3
0046a403
ff868693
02868663
00f00593
0100006f
32075c63
00c42403
00868c63
00442783
ffc7f793
40978733
fee5d4e3
00050613
01092403
00890893
17140863
00442583
00f00713
ffc5f593
409587b3
40f74c63
01192a23
01192823
3e07d663
1ff00793
2eb7ea63
ff85f793
00878793
00492503
00f907b3
0007a683
0055d593
00100713
00b71733
00a76733
ff878593
00b42623
00d42423
00e92223
0087a023
0086a623
40265793
00100593
00f595b3
10b76863
00e5f7b3
02079463
00159593
ffc67613
00e5f7b3
00460613
00079a63
00159593
00e5f7b3
00460613
fe078ae3
00f00813
00361313
00690333
00030513
00c52783
00060e13
2ef50263
0047a703
00078413
00c7a783
ffc77713
409706b3
2ed84263
fe06c2e3
00e40733
00472683
00842603
00098513
0016e693
00d72223
00f62623
00c7a423
11d000ef
00840513
0100006f
00c00793
00f9a023
00000513
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
03010113
00008067
20000693
04000613
03f00513
e65ff06f
00c7a403
00260613
de8794e3
01092403
00890893
e9141ce3
00492703
40265793
00100593
00f595b3
eeb77ce3
00892403
00442b03
ffcb7b13
009b6863
409b07b3
00f00713
14f74663
040077b7
04007cb7
78c7aa83
678ca703
fff00793
01640a33
01548ab3
34f70a63
000017b7
00f78793
00fa8ab3
fffff7b7
00fafab3
000a8593
00098513
044020ef
fff00793
00050b93
28f50c63
29456863
04007c37
750c0c13
000c2583
00ba85b3
00bc2023
00058793
3aaa0463
678ca683
fff00713
3ae68c63
414b8a33
00fa07b3
00fc2023
007bfc93
300c8663
000017b7
419b8bb3
00878593
008b8b93
419585b3
015b8ab3
fff78793
415585b3
00f5fa33
000a0593
00098513
7c9010ef
fff00793
3cf50063
41750533
01450ab3
000c2783
01792423
001aea93
00fa05b3
00bc2023
015ba223
35240863
00f00693
3566f863
00442703
ff4b0793
ff87f793
00177713
00f76733
00e42223
00500613
00f40733
00c72223
00c72423
36f6ee63
004baa83
000b8413
040077b7
7887a703
00b77463
78b7a423
040077b7
7847a703
1ab77663
78b7a223
1a40006f
0014e713
00e42223
009404b3
00992423
0017e793
00098513
00f4a223
714000ef
00840513
e09ff06f
00c42683
00842603
c41ff06f
0095d793
00400713
14f77263
01400713
22f76a63
05c78693
05b78713
00369693
00d906b3
0006a783
ff868693
1cf68863
0047a703
ffc77713
00e5f663
0087a783
fef698e3
00c7a683
00492703
00d42623
00f42423
0086a423
0087a623
cf1ff06f
01400713
12f77663
05400713
1ef76a63
00c4d793
06f78613
06e78513
00361693
c1dff06f
001e0e13
003e7793
00850513
10078e63
00c52783
d09ff06f
00842603
0014e593
00b42223
00f62623
00c7a423
009404b3
00992a23
00992823
0016e793
0114a623
0114a423
00f4a223
00e40733
00098513
00d72023
624000ef
00840513
d19ff06f
0034d613
00848793
b29ff06f
00b405b3
0045a783
00098513
0017e793
00f5a223
5f8000ef
00840513
cedff06f
0014e713
00e42223
009404b3
00992a23
00992823
0017e713
0114a623
0114a423
00e4a223
00b405b3
00098513
00f5a023
5bc000ef
00840513
cb1ff06f
0065d793
03978693
03878713
00369693
ec5ff06f
11240e63
00892403
00442a83
ffcafa93
409a87b3
009ae663
00f00713
e4f748e3
00098513
578000ef
00000513
c6dff06f
05c78613
05b78513
00361693
b01ff06f
00832783
fff60613
1c679263
00367793
ff830313
fe0796e3
00492703
fff5c793
00e7f7b3
00f92223
00159593
c8b7eee3
c8058ce3
00f5f733
00071a63
00159593
00f5f733
004e0e13
fe070ae3
000e0613
b9dff06f
010a8a93
cc1ff06f
00492503
40275593
00100713
00b71733
00a76733
00e92223
e39ff06f
015b85b3
40b005b3
01459593
0145da13
000a0593
00098513
4d5010ef
fff00793
d0f518e3
00000a13
d11ff06f
05400713
08f76263
00c5d793
06f78693
06e78713
00369693
dc5ff06f
15400713
08f76263
00f4d793
07878613
07778513
00361693
a25ff06f
04007c37
750c0c13
000c2783
00fa87b3
00fc2023
c61ff06f
014a1713
c4071ce3
00892403
015b0ab3
001aea93
01542223
cfdff06f
677cac23
c55ff06f
000b8413
cedff06f
00100793
00fba223
eb9ff06f
15400713
06f76263
00f5d793
07878693
07778713
00369693
d3dff06f
55400713
06f76263
0124d793
07d78613
07c78513
00361693
99dff06f
ff8c8c93
019a8ab3
417a8ab3
00000a13
c3dff06f
00840593
00098513
860fc0ef
00892403
000c2583
00442a83
c79ff06f
55400713
02f76463
0125d793
07d78693
07c78713
00369693
cd5ff06f
3f800693
07f00613
07e00513
941ff06f
3f800693
07e00713
cb9ff06f
00492783
e59ff06f
040077b7
1dc7a783
00078067
02058063
04060263
04068863
00064783
00f5a023
00064503
00a03533
00008067
ff010113
00c10593
02060463
02068a63
00064783
00f5a023
00064503
00a03533
01010113
00008067
00000513
00008067
00000513
fedff06f
ffe00513
00008067
ffe00513
fddff06f
00357793
0ff5f693
02078a63
fff60793
02060e63
fff00613
0180006f
00150513
00357713
00070e63
fff78793
02c78063
00054703
fed714e3
00008067
00060793
00300713
02f76663
00079663
00000513
00008067
00f507b3
00c0006f
00150513
fea786e3
00054703
fed71ae3
00008067
0ff5f593
00859713
00b76733
01071893
feff0837
808085b7
00e8e8b3
eff80813
08058593
00300313
00052703
00e8c733
01070633
fff74713
00e67733
00b77733
fa0712e3
ffc78793
00450513
fcf36ee3
f8079ae3
f89ff06f
00b547b3
0037f793
00c508b3
06079663
00300793
06c7f263
00357793
00050713
0c079a63
ffc8f613
40e606b3
02000793
02000293
06d7c263
00058693
00070793
02c77863
0006a803
00478793
00468693
ff07ae23
fec7e8e3
fff60793
40e787b3
ffc7f793
00478793
00f70733
00f585b3
01176863
00008067
00050713
ff157ce3
0005c783
00170713
00158593
fef70fa3
ff1768e3
00008067
0045a683
01c5a783
0005af83
0085af03
00c5ae83
0105ae03
0145a303
0185a803
00d72223
0205a683
01f72023
01e72423
01d72623
01c72823
00672a23
01072c23
00f72e23
02470713
40e607b3
fed72e23
02458593
faf2c6e3
f49ff06f
0005c683
00170713
00377793
fed70fa3
00158593
f0078ee3
0005c683
00170713
00377793
fed70fa3
00158593
fc079ae3
f01ff06f
02a5f663
00c587b3
02f57263
00c50733
0e060a63
fff7c683
fff78793
fff70713
00d70023
fef598e3
00008067
00f00793
02c7e863
00050793
fff60693
0c060c63
00168693
00d786b3
0005c703
00178793
00158593
fee78fa3
fed798e3
00008067
00b567b3
0037f793
0a079063
ff060893
ff08f893
01088893
01150833
00058713
00050793
00072683
01070713
01078793
fed7a823
ff472683
fed7aa23
ff872683
fed7ac23
ffc72683
fed7ae23
fcf81ce3
00c67713
011585b3
00f67813
04070e63
00058713
00078893
00300e13
00072303
00470713
40e806b3
0068a023
00d586b3
00488893
fede64e3
ffc80713
ffc77713
00470713
00367613
00e787b3
00e585b3
f39ff06f
00008067
fff60693
00050793
f31ff06f
00008067
00080613
f1dff06f
00008067
00008067
04c52783
ff010113
00812423
00912223
00112623
01212023
00050413
00058493
02078e63
00249713
00e787b3
0007a503
04050663
00052703
00e7a023
00052823
00052623
00c12083
00812403
00412483
00012903
01010113
00008067
02100613
00400593
295050ef
04a42623
00050793
fa051ae3
00000513
fcdff06f
00100913
00991933
00590613
00261613
00100593
00040513
265050ef
fc050ee3
00952223
01252423
f99ff06f
02058063
0045a703
04c52783
00271713
00e787b3
0007a703
00e5a023
00b7a023
00008067
fd010113
03212023
0105a903
01812423
00010c37
02812423
02912223
01312e23
01412c23
01512a23
01612823
02112623
01712623
00058993
00050a13
00060a93
00068413
01458493
00000b13
fffc0c13
0004ab83
000a8593
00448493
018bf533
ee9f70ef
00850433
000a8593
010bd513
ed9f70ef
01045793
00f50533
01847433
01051793
008787b3
fef4ae23
001b0b13
01055413
fb2b4ee3
02040263
0089a783
04f95863
00490793
00279793
00f987b3
0087a223
00190913
0129a823
02c12083
02812403
02412483
02012903
01812a03
01412a83
01012b03
00c12b83
00812c03
00098513
01c12983
03010113
00008067
0049a583
000a0513
00158593
e39ff0ef
00050493
04050c63
0109a603
00c98593
00c50513
00260613
00261613
bc9ff0ef
0049a703
04ca2783
00271713
00e787b3
0007a703
00e9a023
0137a023
00490793
00048993
00279793
00f987b3
0087a223
00190913
0129a823
f65ff06f
000216b7
00021537
8e068693
00000613
0b500593
96050513
039050ef
fe010113
00812c23
01212823
00058413
00050913
00900593
00868513
00912a23
01312623
01412423
00112e23
01512223
00068493
00060993
00070a13
db9f70ef
00900793
0c97d863
00100793
00000593
00179793
00158593
fea7cce3
00090513
d5dff0ef
00050593
0a050a63
00100793
00f52823
01452a23
00900793
0937d663
00940a93
01340a33
000a8413
00044683
00a00613
00090513
fd068693
dedff0ef
00140413
00050593
ff4412e3
ff898413
008a8433
0299d663
413484b3
009404b3
00044683
00a00613
00090513
fd068693
db9ff0ef
00140413
00050593
fe8492e3
01c12083
01812403
01412483
01012903
00c12983
00812a03
00412a83
00058513
02010113
00008067
00a40413
00900993
fa5ff06f
00000593
f45ff06f
000216b7
00021537
8e068693
00000613
0ce00593
96050513
700050ef
ffff0737
00e57733
00050793
00000513
00071663
01079793
01000513
ff000737
00e7f733
00071663
00850513
00879793
f0000737
00e7f733
00071663
00450513
00479793
c0000737
00e7f733
00071663
00250513
00279793
0007ca63
40000737
00e7f7b3
00150513
00078463
00008067
02000513
00008067
00052783
00050713
0077f693
02068463
0017f693
00000513
04069e63
0027f693
0a068863
0017d793
00f72023
00100513
00008067
01079693
0106d693
00000513
06068e63
0ff7f693
06068063
00f7f693
04068263
0037f693
02068463
0017f693
00069c63
0017d793
00150513
00079663
02000513
00008067
00f72023
00008067
0027d793
0017f693
00250513
fe0696e3
fd5ff06f
0047d793
0037f693
00450513
fa069ee3
fddff06f
0087d793
00f7f693
00850513
fa0690e3
fddff06f
0107d793
0ff7f693
01000513
f80692e3
fddff06f
0027d793
00f72023
00200513
00008067
04c52783
ff010113
00812423
00912223
00112623
00050413
00058493
02078c63
0047a503
06050263
00052703
00e7a223
00c12083
00812403
00100793
00952a23
00052623
00f52823
00412483
01010113
00008067
02100613
00400593
5c8050ef
04a42623
00050793
fa051ce3
000216b7
00021537
8e068693
00000613
14000593
96050513
520050ef
01c00613
00100593
00040513
590050ef
fc050ae3
00100793
00f52223
00200793
00f52423
f85ff06f
fb010113
03312e23
03812423
01062983
0105ac03
04812423
03412c23
04112623
04912223
05212023
03512a23
03612823
03712623
03912223
03a12023
01b12e23
00058a13
00060413
013c4c63
00098713
00058413
000c0993
00060a13
00070c13
00842783
00442583
01898bb3
0177a7b3
00f585b3
a09ff0ef
00a12623
20050a63
00c12783
002b9a93
01478b13
015b0ab3
000b0793
015b7863
0007a023
00478793
ff57ece3
014a0a13
002c1c13
01440793
018a0733
00299993
00f12423
00e12023
013789b3
14ea7863
00400713
01540793
00e12223
1af9f263
000104b7
fff48493
01c0006f
0107dc13
0a0c1063
00012783
004a0a13
004b0b13
10fa7e63
000a2783
0097fd33
fe0d00e3
00812c03
000b0c93
00000413
000c2d83
000ca903
000d0593
009df533
96df70ef
009977b3
00f507b3
000d0593
010dd513
00878433
01095913
951f70ef
01045793
01250533
00f50533
00947433
01051793
0087e7b3
004c0c13
00fca023
004c8c93
01055413
fb3c64e3
00412783
00fb07b3
0087a023
000a2783
0107dc13
f60c04e3
000b2403
00812d83
000b0d13
00040913
00000c93
000da503
000c0593
01095913
00957533
8e5f70ef
012507b3
01978cb3
00947433
010c9613
00866633
00cd2023
002dd503
004d2903
000c0593
8bdf70ef
00997633
010cd793
00c50433
00f40433
004d8d93
004d0d13
01045c93
fb3de4e3
00412783
004a0a13
00fb07b3
0087a023
00012783
004b0b13
eefa66e3
01704863
0180006f
fffb8b93
000b8863
ffcaa783
ffca8a93
fe0788e3
00c12783
04c12083
04812403
0177a823
04412483
04012903
03c12983
03812a03
03412a83
03012b03
02c12b83
02812c03
02412c83
02012d03
01c12d83
00078513
05010113
00008067
408987b3
feb78793
ffc7f793
00478793
00f12223
e4dff06f
000216b7
00021537
8e068693
00000613
15d00593
96050513
24c050ef
fe010113
00812c23
01212823
01312623
00112e23
00912a23
00367793
00060413
00050993
00058913
0a079e63
40245413
06040663
0489a483
0c048a63
00147793
02079063
40145413
04040a63
0004a503
06050663
00050493
00147793
fe0784e3
00048613
00090593
00098513
ce9ff0ef
06090663
00492703
04c9a783
40145413
00271713
00e787b3
0007a703
00e92023
0127a023
00050913
fa041ae3
01c12083
01812403
01412483
00c12983
00090513
01012903
02010113
00008067
00048613
00048593
00098513
c8dff0ef
00a4a023
00052023
00050493
f81ff06f
00050913
f65ff06f
fff78793
00020737
09870713
00279793
00f707b3
0007a603
00000693
f9cff0ef
00050913
f25ff06f
00100593
00098513
ebcff0ef
00050493
02050063
27100793
00f52a23
00100793
00f52823
04a9a423
00052023
f05ff06f
000216b7
00021537
8e068693
00000613
14000593
96050513
0f4050ef
fe010113
01412423
0105aa03
0085a783
01312623
40565993
01498a33
00812c23
00912a23
01212823
01512223
00112e23
001a0913
00058493
00060413
0045a583
00050a93
0127d863
00179793
00158593
ff27cce3
000a8513
e20ff0ef
10050c63
01450813
03305463
00598993
00299993
01350733
00080793
00478793
fe07ae23
fee79ce3
fec98993
01380833
0104a883
01448793
01f47613
00289893
011788b3
0a060463
02000593
40c585b3
00080313
00000693
0007a703
00430313
00478793
00c71733
00d76733
fee32e23
ffc7a683
00b6d6b3
ff17e0e3
01548793
00400713
00f8ea63
409887b3
feb78793
ffc7f793
00478713
00e80833
00d82023
00068463
00090a13
0044a703
04caa783
01c12083
00271713
00e787b3
0007a703
01452823
01812403
00e4a023
0097a023
01012903
01412483
00c12983
00812a03
00412a83
02010113
00008067
0007a703
00478793
00480813
fee82e23
fb17f6e3
0007a703
00478793
00480813
fee82e23
fd17eee3
f95ff06f
000216b7
00021537
8e068693
00000613
1d900593
96050513
765040ef
01052703
0105a783
00050813
40f70533
04f71263
00279793
01480813
01458593
00f80733
00f587b3
0080006f
02e87463
ffc72683
ffc7a603
ffc70713
ffc78793
fec686e3
00c6b6b3
40d006b3
0016e513
00008067
00008067
0105a703
01062783
ff010113
00812423
00912223
01212023
00112623
00058493
00060413
40f70933
1af71463
00279693
01458593
01460713
00d587b3
00d70733
0080006f
18f5fc63
ffc7a603
ffc72683
ffc78793
ffc70713
fed606e3
16d66063
0044a583
c2cff0ef
1a050263
0104ae03
01042583
01448493
002e1e93
01440813
00259593
01450613
000108b7
01252623
01d48eb3
00b805b3
00060f13
00048313
00000f93
fff88893
00032783
00082683
004f0f13
0117f733
01f70733
0116ffb3
41f70733
0106d693
0107d793
40d787b3
41075693
00d787b3
01079693
01177733
00e6e733
00480813
feef2e23
00430313
4107df93
fab86ae3
408586b3
feb68693
01540413
0026d693
00000793
0085e463
00269793
00f607b3
00400813
0085e663
00168693
00269813
010484b3
010608b3
05d4fe63
00010837
00088593
00048613
fff80813
00062783
00458593
00460613
0107f6b3
01f686b3
4106d713
0107d793
00e787b3
01079713
0106f6b3
00d76733
fee5ae23
4107df93
fdd666e3
fffe8e93
409e8eb3
ffcefe93
01d887b3
00071a63
ffc7a703
fffe0e13
ffc78793
fe070ae3
00c12083
00812403
01c52823
00412483
00012903
01010113
00008067
00048793
00100913
00040493
00078413
e95ff06f
fe0946e3
00000913
e89ff06f
00000593
ab0ff0ef
04050263
00c12083
00812403
00100793
00f52823
00052a23
00412483
00012903
01010113
00008067
000216b7
00021537
8e068693
00000613
24000593
96050513
4e5040ef
000216b7
00021537
8e068693
00000613
23200593
96050513
4c9040ef
7ff007b7
00b7f5b3
fcc007b7
00f585b3
00000793
00b05663
00078513
00008067
40b005b3
4145d593
01300793
00b7cc63
000807b7
40b7d5b3
00000793
00078513
00008067
fec58593
01e00713
00100793
00b74663
800007b7
00b7d7b3
00000593
00078513
00008067
fe010113
00912a23
01052483
00812c23
01450413
00249493
009404b3
01212823
ffc4a903
01312623
01412423
00090513
00058993
00112e23
d28ff0ef
02000713
40a707b3
00f9a023
00a00793
ffc48a13
08a7d063
ff550513
05447063
ff84a783
04050063
40a706b3
00d7d733
00a91933
00e96933
ff848613
3ff00737
00e96733
00a797b3
02c47263
ff44a603
00d656b3
00d7e7b3
0140006f
00000793
06051463
3ff00737
00e96733
01c12083
01812403
01412483
01012903
00c12983
00812a03
00078513
00070593
02010113
00008067
00b00693
40a686b3
3ff007b7
00d95733
00f76733
00000793
01447663
ff84a783
00d7d7b3
01550513
00a91933
00f967b3
fa9ff06f
00a91933
3ff00737
00e96733
00000793
f95ff06f
fd010113
01512a23
00058a93
00100593
02912223
01312e23
01412c23
02112623
02812423
03212023
00060493
00068a13
00070993
898ff0ef
10050463
00100737
0144d913
fff70793
7ff97913
00050413
0097f7b3
00090463
00e7e7b3
00f12623
060a9263
00c10513
c58ff0ef
00c12703
00100493
00942823
00e42a23
02050793
08090863
bcd90913
00f90933
03500493
012a2023
40f48533
00a9a023
02c12083
00040513
02812403
02412483
02012903
01c12983
01812a03
01412a83
03010113
00008067
00810513
01512423
bf4ff0ef
00c12703
00050793
04050e63
00812603
02000693
40a686b3
00d716b3
00c6e6b3
00a75733
00d42a23
00e12623
00e034b3
00148493
00e42c23
00942823
f6091ce3
00249713
00e40733
01072503
bce78793
00fa2023
b24ff0ef
00549493
40a48533
f69ff06f
00812683
00d42a23
fc1ff06f
000216b7
00021537
8e068693
00000613
30a00593
96050513
1ed040ef
fd010113
03212023
00058913
00810593
02112623
02812423
02912223
01312e23
00050993
d69ff0ef
00050493
00058413
00090513
00c10593
d55ff0ef
01092703
0109a783
00c12683
40e787b3
00812703
00579793
40d70733
00e787b3
00050713
02f05e63
01479793
00878433
00058693
00048513
00040593
00070613
8f4f50ef
02c12083
02812403
02412483
02012903
01c12983
03010113
00008067
01479793
40f585b3
fc9ff06f
ff010113
01212023
00112623
00812423
00912223
01700793
00050913
04a7da63
00021737
a8072783
a8472583
00021737
a8872403
a8c72483
00078513
00040613
00048693
865f50ef
fff90913
00050793
fe0914e3
00c12083
00812403
00412483
00012903
00078513
01010113
00008067
00020737
00351913
09870713
01270733
01072783
00c12083
00812403
01472583
00412483
00012903
00078513
01010113
00008067
01062683
fff58593
4055d593
00158593
01460793
00269693
00259593
00d786b3
00b505b3
02d7f863
00050713
0007a803
00478793
00470713
ff072e23
fed7e8e3
40c687b3
feb78793
ffc7f793
00478793
00f50533
00b57863
00450513
fe052e23
feb56ce3
00008067
01052703
4055d613
01450693
02c75263
00271713
00e687b3
04f6f263
ffc7a703
ffc78793
fe070ae3
00100513
00008067
00261793
00f687b3
fee650e3
01f5f593
fc058ce3
0007a603
00100513
00b65733
00b71733
fce602e3
00008067
00000513
00008067
fd010113
03212023
02112623
02812423
02912223
01312e23
01412c23
01512a23
01612823
01712623
01812423
00060913
1c058663
00058413
00050993
d15fe0ef
00b90493
01600713
ffc42783
0e977c63
ff84f493
00048713
0e04cc63
0f24ea63
ffc7fa13
ff840a93
12ea5e63
040076b7
26468c13
008c2583
014a8633
00462683
1ec58063
ffe6f593
00b605b3
0045a583
0015f593
14059663
ffc6f693
00da05b3
0ee5d863
0017f793
02079463
ff842b83
417a8bb3
004ba783
ffc7f793
00d786b3
01468b33
36eb5063
00fa0b33
2ceb5263
00090593
00098513
93cfe0ef
00050913
04050c63
ffc42783
ff850713
ffe7f793
00fa87b3
28e78663
ffca0613
02400793
30c7ec63
01300713
22c76063
00050793
00040713
00072683
00d7a023
00472683
00d7a223
00872703
00e7a423
00040593
00098513
8a5fa0ef
00098513
c19fe0ef
01c0006f
01000493
01000713
f124fae3
00c00793
00f9a023
00000913
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00090513
02012903
03010113
00008067
00c62783
00862703
00058a13
00f72623
00e7a423
004aa783
409a06b3
00f00613
0017f793
014a8733
06d66c63
00fa67b3
00faa223
00472783
0017e793
00f72223
00098513
b81fe0ef
00040913
f81ff06f
0017f793
ee0796e3
ff842b83
417a8bb3
004ba783
ffc7f793
ed1ff06f
02812403
02c12083
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00060593
03010113
fe9fd06f
0097e7b3
00faa223
009a85b3
0016e693
00d5a223
00472783
00858593
00098513
0017e793
00f72223
f80fa0ef
f75ff06f
ffc6f693
00da0633
01048593
0eb65063
0017f793
e4079ee3
ff842b83
417a8bb3
004ba783
ffc7f793
00d786b3
01468b33
e2bb4ce3
00cba783
008ba703
ffca0613
02400693
00f72623
00e7a423
008b8913
26c6e063
01300713
00090793
02c77263
00042703
01b00793
00eba423
00442703
00eba623
24c7e663
00840413
010b8793
00042703
00e7a023
00442703
00e7a223
00842703
00e7a423
009b8733
409b07b3
00ec2423
0017e793
00f72223
004ba783
00098513
0017f793
0097e7b3
00fba223
a35fe0ef
e39ff06f
00042683
01b00713
00d52023
00442683
00d52223
18c76663
00840713
00850793
dcdff06f
009a8ab3
409607b3
015c2423
0017e793
00faa223
ffc42783
00098513
00040913
0017f793
0097e7b3
fef42e23
9ddfe0ef
de1ff06f
ffc52783
ffc7f793
00fa0a33
e19ff06f
00cba783
008ba703
ffca0613
02400693
00f72623
00e7a423
008b8913
10c6e063
01300713
00090793
02c77c63
00042703
01b00793
00eba423
00442703
00eba623
10c7fc63
00842783
00fba823
00c42783
00fbaa23
0ad60663
01040413
018b8793
00042703
000b0a13
000b8a93
00e7a023
00442703
00e7a223
00842703
00090413
00e7a423
d91ff06f
00040593
815fe0ef
d0dff06f
00c62783
00862703
02400693
ffca0613
00f72623
00e7a423
008ba703
00cba783
008b8913
00f72623
00e7a423
04c6ee63
01300713
00090793
f8c77ae3
00042703
01b00793
00eba423
00442703
00eba623
06c7fa63
00842703
02400793
00eba823
00c42703
00ebaa23
f4f61ee3
01042703
020b8793
01840413
00ebac23
ffc42703
00ebae23
f49ff06f
00040593
00090513
f7cfe0ef
00090413
000b0a13
000b8a93
ce1ff06f
00842703
00e52423
00c42703
00e52623
00f60e63
01040713
01050793
c31ff06f
00840413
010b8793
f01ff06f
01042683
01840713
01850793
00d52823
01442683
00d52a23
c09ff06f
00040593
00090513
f18fe0ef
dddff06f
00842783
00fba823
00c42783
00fbaa23
00d60863
01040413
018b8793
da5ff06f
01042703
020b8793
01840413
00ebac23
ffc42703
00ebae23
d89ff06f
ff010113
00812423
00912223
00050413
040074b7
00058513
00112623
7804a823
f78f20ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
ff010113
00912223
800004b7
00812423
00112623
fff4c493
00060413
00062023
00b4f6b3
7ff00637
00058793
00050713
06c6d063
00a6e8b3
04088c63
00c5f633
00058813
00000893
02061263
000217b7
a947a683
a907a603
924f50ef
00050713
00058813
00b4f6b3
fca00893
4146d693
801007b7
fff78793
c0268693
00f87833
011686b3
3fe007b7
00f867b3
00d42023
00c12083
00812403
00412483
00070513
00078593
01010113
00008067
f6010113
08c10e93
08f12a23
80000337
ffff07b7
00058e13
fff34313
08d12623
20878793
00810593
000e8693
06112e23
00f12a23
08e12823
09012c23
09112e23
01c12423
01c12c23
00612e23
00612823
01d12223
4c4000ef
00812783
00078023
07c12083
0a010113
00008067
00050e13
04007537
f6010113
67452503
08810e93
08f12a23
80000337
ffff07b7
fff34313
08c12423
08d12623
20878793
00058613
000e8693
00810593
06112e23
00f12a23
08e12823
09012c23
09112e23
01c12423
01c12c23
00612e23
00612823
01d12223
448000ef
00812783
00078023
07c12083
0a010113
00008067
ff010113
00812423
00058413
00e59583
00112623
798040ef
02054063
05042783
00c12083
00a787b3
04f42823
00812403
01010113
00008067
00c45783
fffff737
fff70713
00e7f7b3
00c12083
00f41623
00812403
01010113
00008067
00000513
00008067
00c59783
fe010113
00812c23
00912a23
01212823
01312623
00112e23
1007f713
00058413
00050493
00060913
00068993
04071063
fffff737
fff70713
00e7f7b3
00e41583
00f41623
01812403
01c12083
00098693
00090613
00c12983
01012903
00048513
01412483
02010113
7450306f
00e59583
00200693
00000613
660040ef
00c41783
fb1ff06f
ff010113
00812423
00058413
00e59583
00112623
640040ef
fff00793
02f50463
00c45783
00001737
00c12083
00e7e7b3
04a42823
00f41623
00812403
01010113
00008067
00c45783
fffff737
fff70713
00e7f7b3
00c12083
00f41623
00812403
01010113
00008067
00e59583
1340406f
00b56733
fff00393
00377713
10071063
7f7f87b7
f7f78793
00052603
0005a683
00f672b3
00f66333
00f282b3
0062e2b3
10729263
08d61663
00452603
0045a683
00f672b3
00f66333
00f282b3
0062e2b3
0c729e63
06d61663
00852603
0085a683
00f672b3
00f66333
00f282b3
0062e2b3
0c729863
04d61663
00c52603
00c5a683
00f672b3
00f66333
00f282b3
0062e2b3
0c729263
02d61663
01052603
0105a683
00f672b3
00f66333
00f282b3
0062e2b3
0a729c63
01450513
01458593
f4d60ee3
01061713
01069793
00f71e63
01065713
0106d793
40f70533
0ff57593
02059063
00008067
01075713
0107d793
40f70533
0ff57593
00059463
00008067
0ff77713
0ff7f793
40f70533
00008067
00054603
0005c683
00150513
00158593
00d61463
fe0616e3
40d60533
00008067
00450513
00458593
fcd61ce3
00000513
00008067
00850513
00858593
fcd612e3
00000513
00008067
00c50513
00c58593
fad618e3
00000513
00008067
01050513
01058593
f8d61ee3
00000513
00008067
00b567b3
0037f793
08079263
0005a703
7f7f86b7
f7f68693
00d777b3
00d787b3
00e7e7b3
00d7e7b3
fff00613
06c79e63
00050613
fff00813
00e62023
0045a703
00458593
00460613
00d777b3
00d787b3
00e7e7b3
00d7e7b3
ff0780e3
0005c783
0015c703
0025c683
00f60023
00078a63
00e600a3
00070663
00d60123
00069463
00008067
000601a3
00008067
00050793
0005c703
00178793
00158593
fee78fa3
fe0718e3
00008067
00050613
fb1ff06f
00b567b3
0037f793
00050713
06079863
00300793
06c7f463
feff0337
808088b7
eff30313
08088893
00300e13
0005a683
006687b3
fff6c813
0107f7b3
0117f7b3
02079e63
00d72023
ffc60613
00470713
00458593
fcce6ce3
00158593
00170793
02060463
fff5c683
fff60813
fed78fa3
00068e63
00078713
00080613
00158593
00170793
fe0610e3
00008067
00c70733
00080a63
00178793
fe078fa3
fee79ce3
00008067
00008067
e1010113
1e112623
1f212023
1d812423
1da12023
00058c13
00060913
00d12a23
1e812423
1e912223
1d312e23
1d412c23
1d512a23
1d612823
1d712623
1d912223
1bb12e23
00050d13
ac4fd0ef
00052783
00078513
02f12823
f90f60ef
00cc5783
0e012823
0e012a23
0e012c23
0e012e23
0807f793
02a12623
00078863
010c2783
00079463
3b80106f
10c10793
00078893
0ef12223
000207b7
1c078793
00f12c23
000207b7
3d478793
00090b13
00f12423
000b4783
0e012623
0e012423
02012023
02012a23
02012c23
02012e23
04012223
04012423
00012623
00088c93
22078263
000b0413
02500713
2ce78263
00144783
00140413
fe079ae3
416404b3
21640263
0ec12703
0e812783
016ca023
00970733
00178793
009ca223
0ee12623
0ef12423
00700713
008c8c93
28f74a63
00c12703
00044783
00970733
00e12623
1c078263
fff00313
00144483
0c0103a3
00140413
00000993
00000a13
05a00913
00900a93
02a00b93
00030d93
00140413
fe048793
04f96463
01812703
00279793
00e787b3
0007a783
00078067
00000993
fd048693
00044483
00299793
013787b3
00179793
00f689b3
fd048693
00140413
fedaf2e3
fe048793
fcf970e3
14048463
14910623
0c0103a3
00100a93
00100b93
14c10b13
00012823
00000313
02012423
02012223
00012e23
002a7f93
000f8463
002a8a93
084a7913
0ec12783
00091663
415986b3
40d040e3
0c714703
02070a63
0e812703
0c710693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
2ae6c863
020f8a63
0e812703
0c810693
00dca023
00278793
00200693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
4ce6c2e3
08000713
1ce900e3
41730db3
2bb042e3
100a7713
06071ee3
0e812703
017787b3
016ca023
00170713
017ca223
0ef12623
0ee12423
00700693
36e6cc63
008c8c93
004a7a13
000a0663
415984b3
38904263
0159d463
000a8993
00c12703
01370733
00e12623
300792e3
01012783
0e012423
00078863
01012583
000d0513
b6df90ef
10c10c93
00040b13
000b4783
de0792e3
0ec12783
00078463
2c90106f
00cc5783
0407f793
00078463
32c0206f
1ec12083
1e812403
00c12503
1e412483
1e012903
1dc12983
1d812a03
1d412a83
1d012b03
1cc12b83
1c812c03
1c412c83
1c012d03
1bc12d83
1f010113
00008067
000d0513
fadfc0ef
00452783
00078513
04f12423
c78f60ef
00050793
000d0513
00078493
04f12223
f89fc0ef
00852783
02f12e23
00048463
7b10006f
00044483
dcdff06f
00044483
020a6a13
dc1ff06f
416404b3
d56418e3
00044783
d85ff06f
0e410613
000c0593
000d0513
1d4040ef
f40510e3
10c10c93
d59ff06f
008a7793
000d8313
740790e3
01412783
0b010513
01b12823
00778793
ff87f793
0047a603
0007a583
00878793
00f12a23
6ec090ef
0b012603
0b412683
0b812703
0bc12783
01012303
0f010513
00612823
0ef12e23
0ec12823
0ed12a23
0ee12c23
e55fc0ef
0ca12623
00200793
01012303
00f51463
4780106f
00100793
00f51463
5d80106f
06100793
00f49463
6190106f
04100793
00f49463
0380206f
fdf4f713
fff00793
02e12423
00f31463
1990106f
04700793
00f71463
1a40206f
0fc12d83
05412023
0f012e03
0f412e83
0f812f03
100a6793
000dd463
72d0106f
04012c23
00078a13
00012823
fbf48793
02500713
00f77463
6b40106f
00020737
00279793
32c70713
00e787b3
0007a783
00078067
0e410613
000c0593
000d0513
04612623
05f12023
0a0040ef
0e0516e3
0ec12783
04c12303
04012f83
10c10c93
d29ff06f
0e812483
02012683
00100713
016ca023
00178793
00148493
008c8d93
3ad75ae3
00100713
00eca223
0ef12623
0e912423
00700713
50974ae3
02c12703
03012683
00148493
00e787b3
00eda223
00dda023
0ef12623
0e912423
00700713
008d8d93
509746e3
0f012703
0a010593
0b010513
0ae12823
0f412703
00f12e23
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
6a0060ef
02012783
fff78913
01c12783
360500e3
001b0813
00148493
012787b3
010da023
012da223
0ef12623
0e912423
00700713
008d8d93
30974ae3
03812683
0d410713
00148493
00f687b3
00eda023
00dda223
0ef12623
0e912423
00700713
008d8c93
c8975ae3
0e410613
000c0593
000d0513
771030ef
7a051e63
0ec12783
10c10c93
c75ff06f
01000693
0e812703
0096c463
6d10106f
000206b7
3c468d93
01000913
00700a13
00c0006f
ff048493
04995663
01078793
00170713
01bca023
012ca223
0ef12623
0ee12423
008c8c93
fcea5ee3
0e410613
000c0593
000d0513
705030ef
74051863
ff048493
0ec12783
0e812703
10c10c93
fa994ee3
009787b3
00170713
01bca023
009ca223
0ef12623
0ee12423
00700693
bee6d8e3
0e410613
000c0593
000d0513
6bd030ef
70051463
0ec12783
bd5ff06f
01412783
0c0103a3
0007ab03
00478913
000b1463
25c0106f
fff00793
54fd8ce3
000d8613
00000593
000b0513
01b12a23
fa0fd0ef
00a12823
01412303
00051463
4fd0106f
01012783
41678bb3
0c714783
fffbca93
41fada93
01212a23
00012823
02012423
02012223
00012e23
015bfab3
00000313
a80780e3
001a8a93
a79ff06f
01412703
0c0103a3
00100a93
00072783
00470713
00e12a23
14f10623
00100b93
14c10b13
a3dff06f
01412783
0007a983
00478793
3009dee3
413009b3
00f12a23
00044483
004a6a13
9b1ff06f
01412683
020a7793
00468713
32079ce3
010a7793
00078463
1700106f
040a7793
00078463
3580106f
200a7a13
000a1463
1580106f
01412783
00e12a23
00c12703
0007a783
00040b13
00e78023
af1ff06f
00044483
06c00793
3ef48ee3
010a6a13
94dff06f
01412703
ffff87b7
8307c793
0cf11423
00470793
000d8313
00f12a23
00072d83
000217b7
88c78793
02f12a23
00000913
002a6a93
00200793
07800493
00000693
0cd103a3
fff00693
1cd30863
012de6b3
f7fafa13
1c069063
22031663
04079ee3
001afb93
1b010b13
240b92e3
0c714783
00030a93
01735463
000b8a93
00012823
02012423
02012223
00012e23
ea079ee3
935ff06f
000d8313
010a6a13
020a7793
0c0788e3
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
bffa7a93
00000793
f75ff06f
00044483
06800793
2ef486e3
040a6a13
86dff06f
000d8313
010a6a93
020af793
0a078ae3
01412783
00778b13
ff8b7b13
008b0793
00f12a23
000b2d83
004b2903
00100793
f2dff06f
00044483
008a6a13
82dff06f
00044483
001a6a13
821ff06f
0c714783
00044483
80079ae3
02000793
0cf103a3
809ff06f
00044483
080a6a13
ffcff06f
00044483
00140713
01749463
6190106f
fd048693
00070413
00000d93
fedae063
00044483
002d9793
01b787b3
00179793
00d78db3
fd048693
00140413
fedaf2e3
fbcff06f
02b00793
00044483
0cf103a3
fa8ff06f
000d8313
010a6a13
020a7793
02078ee3
01412783
00778b13
ff8b7b13
004b2783
000b2d83
008b0713
00e12a23
00078913
0407c6e3
fff00793
000a0a93
00f30863
012de7b3
f7fa7a93
6c078263
48091ae3
00900793
49b7e6e3
030d8d93
1bb107a3
000a8a13
00100b93
1af10b13
e5dff06f
000a0a93
00100693
fcd78ae3
00200693
06d78c63
1b010b13
01d91713
007df793
003ddd93
03078793
01b76db3
00395913
fefb0fa3
012de733
000b0613
fffb0b13
fc071ce3
001af693
06068a63
03000693
06d78663
ffe60613
1b010793
fedb0fa3
40c78bb3
000a8a13
00060b13
dedff06f
00100713
00e79463
27d0106f
00200713
000a0a93
f8e798e3
03412683
1b010b13
00fdf793
00f687b3
0007c703
004ddd93
01c91793
01b7edb3
00495913
feeb0fa3
012de7b3
fffb0b13
fc079ce3
1b010793
41678bb3
000a8a13
d91ff06f
06500713
a0975ae3
0f012703
0a010593
0b010513
0ae12823
0f412703
04f12023
0a012023
0ae12a23
0f812703
0a012223
0a012423
0ae12c23
0fc12703
0a012623
0ae12e23
114060ef
04012783
40051663
0e812703
000216b7
8bc68693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
4ce6c6e3
0cc12703
02012683
70d75e63
03012703
02c12683
008c8c93
feecac23
0e812703
00d787b3
fedcae23
00170713
0ef12623
0ee12423
00700693
02e6cae3
02012703
fff70493
ee905463
01000693
0e812703
4896dce3
01000913
00700b93
00c0006f
ff048493
489952e3
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
181030ef
1c051663
0ec12783
0e812703
10c10c93
fb5ff06f
41598933
e5205063
01000613
0e812703
09265463
04812023
01000e13
000c0413
00700d93
00090c13
00030913
00c0006f
ff0c0c13
058e5a63
00812683
01078793
00170713
00dca023
01cca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
00040593
000d0513
101030ef
40051ee3
01000e13
ff0c0c13
0ec12783
0e812703
10c10c93
fb8e4ae3
00090313
000c0913
00040c13
04012403
00812683
012787b3
00170713
00dca023
012ca223
0ef12623
0ee12423
00700693
008c8c93
d8e6d463
0e410613
000c0593
000d0513
04612023
099030ef
0e051263
04012303
0ec12783
10c10c93
41730db3
d7b05263
01000613
0e812703
07b65463
01000313
00700913
00c0006f
ff0d8d93
05b35a63
00812683
01078793
00170713
00dca023
006ca223
0ef12623
0ee12423
008c8c93
fce95ce3
0e410613
000c0593
000d0513
02d030ef
06051c63
01000313
ff0d8d93
0ec12783
0e812703
10c10c93
fbb34ae3
00812683
01b787b3
00170713
00dca023
01bca223
0ef12623
0ee12423
00700693
008c8c93
cce6d663
0e410613
000c0593
000d0513
7d8030ef
02051263
0ec12783
10c10c93
cacff06f
0e410613
000c0593
000d0513
7b8030ef
ce050863
01012583
d0058e63
000d0513
860f90ef
d10ff06f
01000613
0e812703
00d64463
64c0106f
00020637
3c460d93
05212623
04812823
000d8913
000d0413
000a8d93
01000e13
00098a93
00700293
00048993
05f12023
000c0493
00068d13
000b0c13
00030b13
00c0006f
ff0d0d13
05ae5a63
01078793
00170713
012ca023
01cca223
0ef12623
0ee12423
008c8c93
fce2dee3
0e410613
00048593
00040513
714030ef
1a051ae3
01000e13
ff0d0d13
0ec12783
0e812703
10c10c93
00700293
fbae4ae3
000d0693
000b0313
00040d13
000c0b13
04012f83
00048c13
05012403
00098493
000a8993
000d8a93
00090d93
04c12903
00d787b3
00170713
00dca223
01bca023
0ef12623
0ee12423
00700693
008c8c93
b0e6d463
0e410613
000c0593
000d0513
04612623
05f12023
688030ef
ec051ae3
0ec12783
04c12303
04012f83
10c10c93
ad8ff06f
0e410613
000c0593
000d0513
04612023
65c030ef
ea0514e3
0ec12783
04012303
10c10c93
b1cff06f
0cc12603
00c05ae3
01c12703
02012683
00070493
3ee6ce63
02905663
0e812703
009787b3
016ca023
00170713
009ca223
0ef12623
0ee12423
00700693
008c8c93
34e6cee3
fff4c713
41f75713
00e4f4b3
01c12703
409704b3
4c904263
01c12683
400a7713
00db04b3
50071e63
0cc12683
02012703
00e6c663
001a7713
340704e3
03012703
02c12603
008c8c93
feecac23
0e812703
00c787b3
feccae23
00170713
0ef12623
0ee12423
00700613
00e65463
3f00106f
02012703
00eb0833
40d70633
40980933
01265463
00060913
03205863
0e812703
012787b3
009ca023
00170713
012ca223
0ef12623
0ee12423
00700693
008c8c93
00e6d463
4280106f
fff94713
41f75713
00e97933
412604b3
a4905663
01000693
0e812703
7e96de63
01000913
00700b93
00c0006f
ff048493
7e995463
00812683
01078793
00170713
00dca023
012ca223
0ef12623
0ee12423
008c8c93
fcebdce3
0e410613
000c0593
000d0513
4e4030ef
d20518e3
0ec12783
0e812703
10c10c93
fb5ff06f
940316e3
000a8a13
00000313
00000b93
1b010b13
fa8ff06f
001a7613
c4061663
00eca223
0ef12623
0e912423
00700713
ce975a63
0e410613
000c0593
000d0513
48c030ef
cc051ce3
0ec12783
0e812483
10c10d93
cd0ff06f
cd205663
01000713
052758e3
01000b93
00700b13
00c0006f
ff090913
032bdee3
00812703
01078793
00148493
00eda023
017da223
0ef12623
0e912423
008d8d93
fc9b5ce3
0e410613
000c0593
000d0513
424030ef
c60518e3
0ec12783
0e812483
10c10d93
fb5ff06f
01412703
010a7793
00072d83
00470713
00e12a23
14079a63
040a7793
14078263
010d9d93
010ddd93
00000913
f24ff06f
01412703
010af793
00072d83
00470713
00e12a23
02079663
040af793
00078c63
010d9d93
010ddd93
00000913
00100793
e6cff06f
200af793
00078463
0ffdfd93
00000913
00100793
e54ff06f
01412703
010a7793
00072d83
00470713
00e12a23
0c079263
040a7793
0a078a63
010d9d93
410ddd93
41fdd913
00090793
fa07de63
01b037b3
41200933
40f90933
41b00db3
000a0a93
02d00693
00100793
e04ff06f
0e410613
000c0593
000d0513
330030ef
b6051ee3
0ec12783
0e812483
10c10d93
ad0ff06f
0e410613
000c0593
000d0513
30c030ef
b4051ce3
0ec12783
0e812483
10c10d93
ad8ff06f
001a7713
00071463
800ff06f
8ddff06f
000d8313
f10ff06f
00044483
00f12a23
ea1fe06f
03000793
1af107a3
1af10b13
db4ff06f
200a7793
080790e3
41fdd913
00090793
f08ff06f
200a7793
080790e3
00000913
de4ff06f
00c12603
0006a783
00e12a23
41f65693
00c7a023
00d7a223
00040b13
fddfe06f
01412703
00072783
00470713
00e12a23
0007a603
0047a683
0087a703
00c7a783
8e0ff06f
03c12783
00044483
00079463
e19fe06f
0007c783
00079463
e0dfe06f
400a6a13
e05fe06f
00068493
c09044e3
c2dff06f
000d8313
000a0a93
d8cff06f
000217b7
88c78793
000d8313
02f12a23
020a7793
2a078863
01412783
00778b13
ff8b7b13
000b2d83
004b2903
008b0793
00f12a23
001a7793
00078e63
012de7b3
00078a63
03000793
0cf10423
0c9104a3
002a6a13
bffa7a93
00200793
c80ff06f
00144483
200a6a13
00140413
d7dfe06f
0e410613
000c0593
000d0513
1a0030ef
9e0516e3
0ec12783
10c10c93
fb4ff06f
00144483
020a6a13
00140413
d4dfe06f
000217b7
8a078793
000d8313
02f12a23
f61ff06f
000d8313
c84ff06f
04000593
000d0513
a50fc0ef
00ac2023
00ac2823
00051463
3700106f
04000793
00fc2a23
c29fe06f
000b0513
b80f50ef
00050b93
accff06f
01000693
0e812703
5c96dc63
01000b93
00700d93
00c0006f
ff048493
5c9bd263
00812683
01078793
00170713
00dca023
017ca223
0ef12623
0ee12423
008c8c93
fceddce3
0e410613
000c0593
000d0513
0d8030ef
920512e3
0ec12783
0e812703
10c10c93
fb5ff06f
02012703
02412b83
00812e23
00eb0733
05412023
05312623
03512223
02812983
03612423
03c12403
04412a03
04812a83
00700d93
01000913
000c8693
00070b13
080b8663
08099663
fff40413
fffb8b93
0e812703
014787b3
0156a023
00170713
0146a223
0ef12623
0ee12423
00868693
12edcc63
00044603
409b0cb3
01965463
00060c93
03905663
0e812603
019787b3
0096a023
00160613
0196a223
0ef12623
0ec12423
30cdcc63
00044603
00868693
fffcc513
41f55513
00acf733
40e60cb3
01904c63
00c484b3
f60b9ee3
3c0988e3
fff98993
f7dff06f
0e812603
01994863
0580006f
ff0c8c93
05995863
00812703
01078793
00160613
00e6a023
0126a223
0ef12623
0ec12423
00868693
fccddce3
0e410613
000c0593
000d0513
7a5020ef
fe051863
ff0c8c93
0ec12783
0e812603
10c10693
fb994ce3
00812703
019787b3
00160613
00e6a023
0196a223
0ef12623
0ec12423
42cdc0e3
00044603
00868693
00c484b3
f65ff06f
01412703
010a7793
00072d83
00470713
00e12a23
02079263
040a7793
00078a63
010d9d93
010ddd93
00000913
d45ff06f
200a7793
4c079e63
00000913
d35ff06f
0e410613
000c0593
000d0513
70d020ef
f4051c63
0ec12783
10c10693
eb1ff06f
1b010b13
00000793
00812823
00912e23
000b0413
03312223
000c0b13
000d8493
00090993
03c12d83
400afa13
0ff00b93
00030c13
00078913
0240006f
00a00613
00000693
00048513
00098593
2d9040ef
3e098463
00050493
00058993
00a00613
00000693
00048513
00098593
078050ef
03050513
fea40fa3
00190913
fff40413
fa0a0ee3
000dc683
fad91ae3
fb7908e3
36099463
00900793
3697e063
000c0313
1b010793
000b0c13
00040b13
01c12483
02412983
01012403
03b12e23
03212023
41678bb3
000a8a13
920ff06f
0e812703
000216b7
8bc68693
00dca023
00178793
00100693
00170713
00dca223
0ef12623
0ee12423
00700693
008c8c93
06e6ce63
1e061863
02012683
001a7713
00d76733
00071463
af9fe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
60e6c263
02012683
00170713
0168a023
00f687b3
00d8a223
0ef12623
0ee12423
00700693
00888c93
00e6c463
a9dfe06f
e09fe06f
0e410613
000c0593
000d0513
575020ef
dc051063
0cc12603
0ec12783
10c10c93
f69ff06f
00040d13
00048c13
da4ff06f
0e410613
000c0593
000d0513
545020ef
d8051863
0ec12783
10c10c93
b1cff06f
00812683
009787b3
009ca223
00dca023
00170713
0ef12623
0ee12423
00700693
00e6c463
a1dfe06f
d8dfe06f
0e410613
000c0593
000d0513
4f9020ef
d4051263
00044603
0ec12783
10c10693
cd5ff06f
00040c13
d2cff06f
0f012783
0a010593
0b010513
0af12823
0f412783
0a012023
0a012223
0af12a23
0f812783
0a012423
0a012623
0af12c23
0fc12783
0af12e23
56c050ef
320540e3
0c714783
04700713
1c975e63
00021837
88080b13
00012823
02012423
02012223
00012e23
f7fa7a13
00300a93
00300b93
00000313
00078463
e2dfe06f
8a5fe06f
01412783
00040b13
0007a783
00e12a23
00c12703
00e7a023
99dfe06f
00600793
000d8b93
1bb7e663
00021837
000b8a93
01212a23
8b480b13
855fe06f
00812703
012787b3
00148493
00eda023
c4dfe06f
03012703
02c12683
008c8893
00eca023
0e812703
00f687b3
00dca223
00170713
0ef12623
0ee12423
00700693
42e6c663
e20654e3
ff000693
40c004b3
3ed658e3
01000913
00700b93
00c0006f
ff048493
3c995ee3
00812683
01078793
00170713
00d8a023
0128a223
0ef12623
0ee12423
00888893
fcebdce3
0e410613
000c0593
000d0513
385020ef
bc051863
0ec12783
0e812703
10c10893
fb5ff06f
0fc12783
3a07d863
02d00793
0cf103a3
04700713
229750e3
00021837
88880b13
ec9ff06f
00812683
009787b3
00170713
00dca023
009ca223
0ef12623
0ee12423
00700693
008c8c93
d2e6de63
0e410613
000c0593
000d0513
315020ef
b6051063
0ec12783
10c10c93
d1cff06f
04412783
04812583
00000913
40f40433
00078613
00040513
ca4fe0ef
001dc583
00a00613
00000693
00b03833
00048513
00098593
010d8db3
6f4040ef
c21ff06f
00900793
c097ece3
c5dff06f
00021837
87c80b13
e29ff06f
0e410613
000c0593
000d0513
29d020ef
ae051463
0ec12783
10c10c93
c8cff06f
00600b93
e55ff06f
02012703
00eb0833
40d70633
40980933
d3265463
00060913
d20ff06f
01412783
00e12a23
00c12703
0007a783
00040b13
00e79023
fa8fe06f
0ffdfd93
00000913
859ff06f
018d9d93
418ddd93
41fdd913
00090793
e85fe06f
0ffdfd93
00000913
d65fe06f
00030693
00200613
0b010a93
0d010793
0cc10713
0dc10813
000a8593
000d0513
04612823
04d12623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
0bb12e23
c30fa0ef
02812703
04700793
01c12f03
02012e83
02412e03
04c12683
05012303
00050b13
64f70863
04600793
00d50933
06f71ee3
00054703
03000793
2ef700e3
0a010b93
0cc12783
00f90933
000b8593
000a8513
00612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
0a012023
0a012223
0a012423
0a012623
01c050ef
01c12303
00090693
02050263
0dc12683
0126fe63
03000713
00168793
0cf12e23
00e68023
0dc12683
ff26e8e3
416687b3
02f12023
0cc12703
04700793
00e12e23
02812703
52f70463
02812703
04600793
02f700e3
01c12783
02812603
04100693
fff78b93
0d712623
0ff4f793
00000713
00d61863
00f78793
0ff7f793
00100713
0cf10a23
02b00793
000bda63
01c12783
00100b93
40fb8bb3
02d00793
0cf10aa3
00900793
0b77d6e3
0e310a13
000a0913
00a00593
000b8513
d9cf40ef
03050793
fef90fa3
000b8513
00a00593
d04f40ef
000b8a93
06300793
00090d93
00050b93
fff90913
fd57c6e3
03050693
0ff6f693
ffed8793
fed90fa3
2947f0e3
0d610713
0080006f
0007c683
00d70023
00178793
00170713
ff4798e3
0e510793
0d610713
41b787b3
00f707b3
0d410713
40e787b3
02f12c23
02012703
03812683
00100793
00d70bb3
0ce7d6e3
02c12783
00fb8bb3
04012783
fffbca93
41fada93
bff7fa13
100a6a13
015bfab3
02012423
02012223
00012e23
05812783
40078a63
02d00793
0cf103a3
00000313
001a8a93
c18fe06f
0e410613
000c0593
000d0513
7c0020ef
d2cfe06f
0c714783
c59ff06f
0e410613
000c0593
000d0513
7a4020ef
00050463
fedfe06f
0cc12603
0ec12783
0e812703
10c10893
9c065ce3
bb1ff06f
00600313
e74fe06f
00130693
00200613
d5dff06f
00030693
00300613
d51ff06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
695070ef
0cc10613
bddfd0ef
00058613
00050593
000a8513
485070ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
0e8050ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
549040ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000217b7
8a078793
02f12223
fff30913
06912023
07312423
07912823
07a12a23
07812c23
01c12483
00090c13
04812e23
07412223
06612623
000b0c93
07612e23
00068d13
000e0d93
000e8913
000f0993
0480006f
000b8593
000a8513
02c12023
01f12e23
0bf12c23
0ac12e23
0b612823
0b412a23
0a012023
0a012223
0a012423
0a012623
4a1040ef
fffc0c13
00090f93
00098613
0e050263
400307b7
00048613
000b8593
000a8513
08f12e23
0ba12023
0bb12223
0b212423
0b312623
08012823
08012a23
08012c23
7b1040ef
000a8513
089070ef
00050593
00050413
000a8513
0b012a03
0b412983
0b812b03
0bc12903
17d070ef
0b012683
04c12603
00048593
08d12023
0b412683
000b8513
09412823
08d12223
0b812683
09312a23
09612c23
08d12423
0bc12683
09212e23
08d12623
30c060ef
02412783
0a012b03
0a412a03
008786b3
0006c683
0a812f83
0ac12603
05912a23
00dc8023
05812823
fff00793
001c8c93
000b0d13
000a0d93
000f8913
00060993
eefc10e3
06c12303
000b0393
000a0293
3ffe0937
000b8593
000a8513
02612023
00812e23
06012483
05c12403
06412a03
0a712823
06712223
0a512a23
06512023
0bf12c23
05f12e23
0ac12e23
04c12623
0a012023
0a012223
0a012423
0b212623
41d040ef
000c8d93
06812983
07012c83
07412d03
07812c03
07c12b03
02012303
40a04463
000b8593
000a8513
325040ef
02012303
00051863
01c12783
0017f913
3e091463
05012783
03000693
00178713
00ed8733
0007c863
001d8d93
fedd8fa3
ffb71ce3
416d87b3
02f12023
b01ff06f
02812b03
02012703
02812e23
04012a03
00eb0733
01c12403
04c12983
02412a83
00068c93
00976463
e25fe06f
00070493
e1dfe06f
01c12703
ffd00793
00f74463
02e35463
ffe48493
fdf4f793
02f12423
acdff06f
0c714783
00000313
00078463
d90fe06f
808fe06f
02012783
01c12703
30f74263
04012783
01c12703
0017f793
00070b93
00078663
02c12783
00f70bb3
04012783
4007f793
00078663
01c12783
44f04463
fffbca93
41fada93
015bfab3
06700493
02012423
02012223
b81ff06f
04012783
00d50933
0017f793
22079663
0dc12683
a21ff06f
0e410613
000c0593
000d0513
340020ef
00050463
b89fe06f
00044603
0ec12783
10c10693
00c484b3
b2cff06f
07800793
03000713
0ce10423
002a6713
0cf104a3
04e12023
06300793
00012823
14c10b13
3667c863
0fc12d83
fdf4f793
02f12423
04012c23
0f012e03
0f412e83
0f812f03
102a6a13
120dc063
06100793
00f48463
9f0fe06f
0b010a93
000a8513
04612e23
0bc12823
0bd12a23
0be12c23
0bb12e23
1fd070ef
0cc10613
f44fd0ef
00058613
00050593
000a8513
7ec070ef
09010793
00078593
00f12e23
0b012783
0a010b93
08010613
08f12823
0b412783
000b8513
04c12623
08f12a23
0b812783
08012023
08012223
08f12c23
0bc12783
08012423
08f12e23
3ffc07b7
08f12623
451040ef
0a012683
0a412e03
0a812e83
0ac12f03
000b8593
000a8513
0ad12823
04d12a23
0bc12a23
05c12823
0bd12c23
03d12223
0be12e23
03e12023
0a012023
0a012223
0a012423
0a012623
0b1040ef
02012f03
02412e83
05012e03
05412683
05c12303
00051663
00100793
0cf12623
000217b7
88c78793
02f12223
b69ff06f
00012823
00078a13
800007b7
01b7cdb3
02d00793
04f12c23
ed5ff06f
0e410613
000c0593
000d0513
198020ef
00050463
9e1fe06f
0cc12683
0ec12783
10c10c93
bf1fe06f
02d00793
0cf103a3
ce0ff06f
0c714783
01212a23
02012423
02012223
00012e23
00030a93
00030b93
00000313
00078463
b18fe06f
d91fd06f
00020637
3c460d93
a7dfe06f
00021837
88480b13
cacff06f
0a010b93
f9cff06f
0e410613
000c0593
000d0513
118020ef
00050463
961fe06f
0cc12483
02012703
0ec12783
10c10c93
40970633
bb1fe06f
05800793
dd5ff06f
04012783
01c12703
0017f793
0067e7b3
2ae05063
28079463
01c12b83
06600493
04012783
4007f793
18079663
fffbca93
41fada93
015bfab3
d45ff06f
02012783
02c12703
06700493
00e78bb3
01c12783
fcf048e3
40fb8bb3
001b8b93
fffbca93
41fada93
015bfab3
d15ff06f
000206b7
3c468d93
990fe06f
000a0a93
cf0fe06f
05412783
000d8713
0cf12e23
02412783
fffdc683
00f7c603
02d61063
03000593
feb70fa3
0dc12703
fff70793
0cf12e23
fff74683
fed606e3
00168613
03900593
0ff67613
00b68663
fec70fa3
bf1ff06f
02412783
00a7c603
fec70fa3
be1ff06f
0d610793
00071863
03000793
0cf10b23
0d710793
1b010713
030b8b93
40e78733
01778023
0dd70793
02f12c23
fb8ff06f
00812683
009787b3
00170713
00d8a023
0098a223
0ef12623
0ee12423
00700693
00888893
a0e6d463
0e410613
000c0593
000d0513
7a9010ef
00050463
ff0fe06f
0ec12783
0e812703
10c10893
9e0ff06f
00130593
000d0513
00612823
878fb0ef
01012303
00050b13
1a050e63
00a12823
c75ff06f
00030463
e5dfd06f
00100313
e55fd06f
fff00793
00f12623
cd1fd06f
04012783
0017f793
f2078c63
f2cff06f
06700493
03c12603
0ff00713
00064783
16e78463
01c12683
00000513
00000593
00d7de63
40f686b3
00164783
04078463
00158593
00160613
fee794e3
02c12e23
00d12e23
02b12223
02a12423
02812783
02412703
04412583
00e78533
b31f30ef
01750bb3
fffbca93
41fada93
015bfab3
ee4ff06f
00064783
00150513
fbdff06f
0a010b93
000b8593
000a8513
04612623
0bc12823
03c12223
0bd12a23
03d12023
0be12c23
01e12e23
04d12823
0bb12e23
0a012023
0a012223
0a012423
0a012623
538040ef
01c12f03
02012e83
02412e03
04c12303
cc050a63
05012683
00100793
40d787b3
0cf12623
cc4ff06f
02c12783
06600493
00f70bb3
006b8bb3
d75ff06f
00079a63
00100a93
06600493
00100b93
abdff06f
02c12783
06600493
00178b93
006b8bb3
fffbca93
41fada93
015bfab3
a9dff06f
01412783
0007ad83
00478793
000dd463
fff00d93
00144483
00f12a23
00070413
9b5fd06f
00200793
02f12c23
db4ff06f
00c00793
00fd2023
fff00793
00f12623
b49fd06f
02012423
02012223
ecdff06f
00cc5783
0407e793
00fc1623
b1dfd06f
0645a703
fd010113
000027b7
01612823
02112623
02812423
02912223
03212023
01312e23
01412c23
01512a23
01712623
01812423
00e7f7b3
00060b13
0a078863
00862783
00062b83
00058913
00050993
fff00a93
08078863
004bac03
000ba403
002c5a13
060a0663
00000493
00c0006f
00440413
049a0c63
00042583
00090613
00098513
125010ef
00148493
ff5512e3
fff00513
02c12083
02812403
000b2423
000b2223
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
008b2783
ffcc7c13
418787b3
00fb2423
008b8b93
f6079ce3
00000513
fadff06f
88df70ef
fa5ff06f
00862703
00070463
f05ff06f
00062223
00000513
00008067
ed010113
11312e23
11512a23
11712623
12112623
12812423
12912223
13212023
11412c23
11612823
11812423
11912223
11a12023
0fb12e23
00d12823
00050a93
00058993
00060b93
00050663
03852783
62078663
00c99703
000026b7
01071793
0107d793
00d7f633
02061863
0649a603
00d767b3
01079793
ffffe737
4107d793
fff70713
00e67733
00f99623
01079793
06e9a223
0107d793
0087f713
3e070a63
0109a703
3e070663
01a7f793
00a00713
40e78063
000207b7
3e478793
00020b37
04c10493
00f12a23
00020937
550b0793
000b8c13
04912023
04012423
04012223
00012c23
00012e23
02012223
02012023
00012623
00f12423
56090913
00048b93
000c4783
26078263
000c0413
02500713
46e78263
00144783
00140413
fe079ae3
41840cb3
25840263
04812703
04412783
018ba023
00ec8733
00178793
019ba223
04e12423
04f12223
00700693
008b8b93
02f6d063
420700e3
04010613
00098593
000a8513
d91ff0ef
20051463
00048b93
00c12703
00044783
01970733
00e12623
1e078463
00144683
00140c13
02010da3
fff00a13
00012223
00000b13
05a00c93
00900d13
02a00613
001c0c13
fe068793
04fce863
01412703
00279793
00e787b3
0007a783
00078067
00012223
fd068793
00412583
000c4683
001c0c13
00259713
00b70733
00171713
00e787b3
00f12223
fd068793
fcfd7ee3
fe068793
fafcfce3
16068463
08d10623
02010da3
00100c93
00100d13
08c10413
00000a13
002b7f93
000f8463
002c8c93
04412703
084b7f13
04812783
00170693
00068613
000f1863
00412583
41958db3
0fb04ce3
03b14683
02068a63
03b10713
00178793
00eba023
00100713
00eba223
04f12423
04c12223
00700713
04c748e3
00060713
008b8b93
00160613
040f8c63
03c10713
00278793
00eba023
00200713
00eba223
04f12423
04c12223
00700713
08c750e3
32078ce3
04010613
00098593
000a8513
03e12423
c35ff0ef
0a051663
04412703
04812783
02812f03
00048b93
00170613
08000693
62df0a63
41aa0a33
71404263
00fd07b3
008ba023
01aba223
04f12423
04c12223
00700713
60c75463
12078ee3
04010613
00098593
000a8513
bddff0ef
04051a63
04812783
00048b93
004b7e13
000e0863
00412703
41970d33
13a044e3
00412403
01945463
000c8413
00c12703
00870733
00e12623
74079463
000c4783
04012223
00048b93
da0792e3
04812783
5e079ae3
00c9d783
0407f793
620792e3
12c12083
12812403
00c12503
12412483
12012903
11c12983
11812a03
11412a83
11012b03
10c12b83
10812c03
10412c83
10012d03
0fc12d83
13010113
00008067
000a8513
e4cfa0ef
00452783
00078513
02f12023
b19f30ef
00050793
000a8513
00078413
02f12223
e28fa0ef
00852783
02a00613
00f12e23
320416e3
000c4683
dadff06f
000c4683
020b6b13
da1ff06f
010b6b13
020b7793
1a078063
01012783
00778793
ff87f793
0047a683
0007ad03
00878793
00f12823
00068c93
1a06c863
fff00693
000b0d93
00da0863
019d66b3
f7fb7d93
120688e3
1a0c9ae3
00900693
1ba6e6e3
030d0793
0ef107a3
000d8b13
00100d13
0ef10413
000a0c93
01aa5463
000d0c93
03b14783
00f037b3
00fc8cb3
d91ff06f
00098593
000a8513
da8f60ef
500510e3
00c9d783
00a00713
01a7f793
c0e794e3
00e99783
c007c0e3
12812403
01012683
12c12083
12412483
12012903
11812a03
11012b03
10812c03
10412c83
10012d03
0fc12d83
000b8613
00098593
10c12b83
11c12983
000a8513
11412a83
13010113
4e90006f
010b6b13
020b7793
06078c63
01012783
00778793
ff87f793
0007ad03
0047ac83
00878793
00f12823
bffb7d93
00000693
00000613
02c10da3
fff00613
0cca0863
019d6633
f7fdfb13
5e061663
340a1463
02069ae3
001dfd13
0f010413
f00d0ae3
03000793
0ef107a3
0ef10413
f05ff06f
41840cb3
bb8418e3
00044783
c01ff06f
01012683
010b7713
0006a783
00468693
00d12823
14071e63
040b7713
14070663
01079d13
010d5d13
00000c93
f7dff06f
01012683
010b7713
0006a783
00468693
00d12823
14071063
040b7713
12070863
01079d13
410d5d13
41fd5c93
000c8693
e406dce3
02d00613
01a036b3
41900733
02c10da3
fff00613
40d70cb3
41a00d33
000b0d93
00100693
f2ca1ce3
00100613
e4c680e3
00200613
28c68863
0f010413
01dc9793
007d7693
003d5d13
03068693
01a7ed33
003cdc93
fed40fa3
019d67b3
00040593
fff40413
fc079ce3
001df793
28078663
03000793
28f68263
ffe58593
fef40fa3
0f010793
40b78d33
000d8b13
00058413
dfdff06f
d01f60ef
9d5ff06f
01012783
02010da3
0007a403
00478d93
20040ce3
fff00793
16fa02e3
000a0613
00000593
00040513
f15fa0ef
2c0502e3
40850d33
01b12823
00000a13
db5ff06f
01012703
02010da3
00100c93
00072783
00470713
00e12823
08f10623
00100d13
08c10413
b31ff06f
200b7713
24071ae3
00078d13
00000c93
e31ff06f
200b7713
220710e3
41f7dc93
00078d13
000c8693
d25ff06f
01012783
0007a703
00478793
00e12223
78075463
00412703
00f12823
40e00733
00e12223
000c4683
004b6b13
a65ff06f
000c4683
06c00793
12f68ae3
010b6b13
a51ff06f
000c4683
06800793
10f688e3
040b6b13
a3dff06f
010b6d93
020df793
62078063
01012783
00100693
00778793
ff87f793
0007ad03
0047ac83
00878793
00f12823
d99ff06f
000c4683
001b6b13
a01ff06f
03b14783
000c4683
9e079ae3
02000793
02f10da3
9e9ff06f
000c4683
080b6b13
9ddff06f
000c4683
001c0713
1cc688e3
fd068793
00070c13
00000a13
9cfd62e3
000c4683
002a1713
01470a33
001a1a13
00fa0a33
fd068793
001c0c13
fefd72e3
9a1ff06f
02b00793
000c4683
02f10da3
98dff06f
01012783
ffff86b7
8306c693
0007ad03
00478793
00f12823
000217b7
88c78793
02d11e23
00000c93
002b6d93
00f12c23
00200693
ce1ff06f
01012683
020b7793
00468713
6a079063
010b7793
020794e3
040b7793
08079ce3
200b7e13
000e0ce3
01012783
00e12823
00c12703
0007a783
00e78023
86dff06f
00100613
0ec68ce3
00200613
000b0d93
d6c69ce3
01812683
0f010413
00fd7793
00f687b3
0007c703
004d5d13
01cc9793
01a7ed33
004cdc93
fee40fa3
019d67b3
fff40413
fc079ce3
0f010793
40878d33
000d8b13
b89ff06f
00100713
000d0793
04812623
05a12823
05a12423
04e12223
00048b93
008b8b93
a19ff06f
00412683
41968db3
9db054e3
01000693
07b6dc63
01000e93
00700f13
0180006f
00270613
008b8b93
00068713
ff0d8d93
05bedc63
01078793
00170693
012ba023
01dba223
04f12423
04d12223
fcdf5ae3
14078863
04010613
00098593
000a8513
d80ff0ef
9e051ce3
04412703
01000e93
ff0d8d93
04812783
00048b93
00170613
00700f13
fbbec8e3
01b787b3
012ba023
01bba223
04f12423
04c12223
00700713
00060593
52c75e63
70078e63
04010613
00098593
000a8513
d28ff0ef
9a0510e3
04412703
41aa0a33
04812783
00048b93
00170613
914052e3
01000693
0746da63
01000893
00700d93
0180006f
00270613
008b8b93
00068713
ff0a0a13
0548da63
01078793
00170693
012ba023
011ba223
04f12423
04d12223
fcdddae3
04078e63
04010613
00098593
000a8513
cb4ff0ef
920516e3
04412703
01000893
ff0a0a13
04812783
00048b93
00170613
fb48cae3
014787b3
012ba023
014ba223
04f12423
04c12223
00700713
2cc74663
008b8b93
00160613
865ff06f
00100613
00000713
00048b93
f75ff06f
04010613
00098593
000a8513
c4cff0ef
8a0506e3
8c1ff06f
00100613
00000713
00048b93
e81ff06f
32078863
04010613
00098593
000a8513
03e12623
03f12423
c18ff0ef
880518e3
04412703
04812783
02c12f03
02812f83
00048b93
00170613
f88ff06f
3a079e63
03b14703
5e071463
2e0f8663
03c10793
04f12623
00200793
04f12823
00100613
00048b93
00060713
008b8b93
00170613
fa8ff06f
000b0d93
ad5ff06f
01000613
65b65063
000b8613
01000e93
00040b93
00700293
00098413
03f12423
000d8993
000c0d93
000a0c13
000f0a13
01c0006f
00270513
00860613
00068713
ff098993
053ede63
00170693
00812583
01078793
01d62223
00b62023
04f12423
04d12223
fcd2d8e3
08078663
04010613
00040593
000a8513
b3cff0ef
4a051863
04412703
01000e93
ff098993
04812783
00048613
00170513
00700293
fb3ec6e3
02812f83
000a0f13
00050593
000c0a13
000d8c13
00098d93
00040993
000b8413
00060b93
00812703
01b787b3
01bba223
00eba023
04f12423
04b12223
00700713
eeb740e3
008b8b93
00158613
00058713
e1cff06f
00000713
00100513
00048613
f41ff06f
04012223
004b7e13
0e0e0063
00412703
41970d33
0da05a63
00048b93
01000713
04412683
53a75263
01000d93
00700413
0180006f
00268613
008b8b93
00070693
ff0d0d13
05adda63
00812603
01078793
00168713
00cba023
01bba223
04f12423
04e12223
fce458e3
06078863
04010613
00098593
000a8513
a38ff0ef
ea051863
04412683
ff0d0d13
04812783
00048b93
00168613
fbadcae3
00812703
01a787b3
01aba223
00eba023
04f12423
04c12223
00700713
e4c75263
02078863
04010613
00098593
000a8513
9e8ff0ef
e6051063
04812783
e24ff06f
00100613
00000693
00048b93
f5dff06f
00412403
01945463
000c8413
00c12783
008787b3
00f12623
e14ff06f
ba0784e3
04010613
00098593
000a8513
99cff0ef
e0051a63
04412603
04812783
00048b93
00160613
d7cff06f
04012223
00048b93
bf4ff06f
ee0a1063
000d8b13
00000a13
00000d13
0f010413
ee0ff06f
01012683
010df713
0006a783
00468693
00d12823
02071463
040df713
00070c63
01079d13
010d5d13
00000c93
00100693
f6cff06f
200df713
38071063
00078d13
00000c93
00100693
f54ff06f
00100613
00000713
00048b93
cecff06f
140f9463
00000713
00100613
00048b93
cd8ff06f
400df793
03412423
03312623
000c8a13
000d0993
00000b13
01c12d03
0f010413
00078c93
0240006f
00a00613
00000693
00098513
000a0593
289020ef
280a0463
00050993
00058a13
00a00613
00000693
00098513
000a0593
028030ef
03050513
fea40fa3
001b0b13
fff40413
fa0c8ee3
000d4683
fb669ae3
0ff00793
fafb06e3
180a1863
00900793
1937e463
0f010793
01a12e23
02812a03
02c12983
40878d33
000d8b13
dc8ff06f
000c4683
00f12823
af0ff06f
04010613
00098593
000a8513
03e12623
03f12423
824ff0ef
c8051e63
04412703
04812783
02c12f03
02812f83
00048b93
00170613
b5cff06f
008b8b93
00160613
00058713
be4ff06f
00c12603
0006a783
00e12823
41f65693
00c7a023
00d7a223
9e4ff06f
01c12783
000c4683
a8078063
0007c783
a6078c63
400b6b13
a70ff06f
03c10793
04f12623
00200793
04f12823
00100713
00048b93
bd9ff06f
000b0d93
819ff06f
000217b7
88c78793
00f12c23
020b7793
06078063
01012783
00778793
ff87f793
0007ad03
0047ac83
00878793
00f12823
001b7613
00060e63
019d6633
00060a63
03000613
02c10e23
02d10ea3
002b6b13
bffb7d93
00200693
d7cff06f
000217b7
8a078793
00f12c23
020b7793
fa0794e3
01012603
010b7713
00062783
00460613
00c12823
06071e63
040b7713
06070663
01079d13
010d5d13
00000c93
f95ff06f
00040513
ee5f20ef
00050d13
01b12823
00000a13
c60ff06f
02412783
02012583
00000b13
40f40433
00078613
00040513
e28fc0ef
001d4583
00a00613
00000693
00b03733
00098513
000a0593
00ed0d33
079020ef
df5ff06f
200b7713
0c071e63
00078d13
00000c93
f29ff06f
00040993
b00ff06f
001c4683
200b6b13
001c0c13
928ff06f
001c4683
020b6b13
001c0c13
918ff06f
01012783
0007a783
00e12823
00c12703
00e7a023
858ff06f
00600793
000a0d13
0347ea63
00021337
000d0c93
01b12823
8b430413
950ff06f
00900793
d737ece3
dc1ff06f
00100613
00000713
00048b93
a00ff06f
00600d13
fcdff06f
03b10793
04f12623
00100793
04f12823
00100613
00048b93
970ff06f
01012783
00e12823
00c12703
0007a783
00e79023
fe1fe06f
01879d13
418d5d13
41fd5c93
000c8693
b04ff06f
0ff7fd13
00000c93
e51ff06f
0ff7fd13
00000c93
be0ff06f
0ff7fd13
00000c93
00100693
bd8ff06f
04010613
00098593
000a8513
d89fe0ef
a00ff06f
000a0d13
01b12823
00000a13
af4ff06f
00068593
a7dff06f
00168613
b4dff06f
000b0d93
ac8ff06f
fff00793
00f12623
9d8ff06f
01012783
0007aa03
00478793
000a5463
fff00a13
001c4683
00f12823
00070c13
fe1fe06f
04007737
00050793
67472503
00060693
00058613
00078593
e1dfe06f
00c5d783
0645ae03
00e5d303
01c5a883
0245a803
b8010113
ffd7f793
40000713
46812c23
00f11a23
00058413
07010793
00810593
46912a23
47212823
46112e23
00050913
07c12623
00611b23
03112223
03012623
00f12423
00f12c23
00e12823
00e12e23
02012023
db1fe0ef
00050493
02055c63
01415783
0407f793
00078863
00c45783
0407e793
00f41623
47c12083
47812403
47012903
00048513
47412483
48010113
00008067
00810593
00090513
c9df50ef
fc0500e3
fff00493
fb9ff06f
040077b7
1d87a783
00078067
02058463
0ff00793
00c7e863
00c58023
00100513
00008067
08a00793
00f52023
fff00513
00008067
00000513
00008067
ff010113
00058713
00812423
00912223
00060593
00050413
040074b7
00068613
00070513
00112623
7804a823
f3cee0ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
040077b7
6747a703
ff010113
00068793
00060813
00112623
00c72883
00050693
00058713
00078613
02080063
000217b7
9b478793
000215b7
9c458593
00088513
390000ef
45d010ef
00020837
70c80793
70c80813
fe1ff06f
ff010113
00060693
00000613
00112623
f99ff0ef
00050593
00000693
00000613
00000513
43d0106f
fe010113
00812c23
00112e23
00912a23
01212823
01312623
0105d693
00058793
00050413
01065713
0c069c63
12071863
01061593
01079513
0105d593
01055513
cdcf20ef
00050593
00040513
979f90ef
00050413
04050863
ffc52603
02400713
ffc67613
ffc60613
04c76e63
01300693
00050793
02c6f263
00052023
00052223
01b00793
06c7f463
00052423
00052623
01050793
0ce60a63
0007a023
0007a223
0007a423
01c12083
00040513
01812403
01412483
01012903
00c12983
02010113
00008067
00000593
ea8f20ef
01c12083
00040513
01812403
01412483
01012903
00c12983
02010113
00008067
00850793
0007a023
0007a223
0007a423
fa9ff06f
06071c63
00068913
00060993
01079513
01061593
0105d593
01055513
c00f20ef
00050493
01091593
01099513
0105d593
01055513
be8f20ef
0104d793
00f505b3
0105d793
02079a63
01049493
01059593
0104d493
0095e5b3
ef1ff06f
00070913
00058993
fa9ff06f
00052823
01850793
00052a23
f25ff06f
074000ef
00c00793
00f52023
00000413
f1dff06f
ff010113
00812423
00912223
00050413
040074b7
00058513
00112623
7804a823
124020ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
040077b7
6747a503
00008067
ff010113
00112623
00812423
00912223
01212023
02058063
00058413
00050493
00050663
03852783
0a078c63
00c41783
02079263
00c12083
00812403
00000913
00412483
00090513
00012903
01010113
00008067
00040593
00048513
eacf50ef
02c42783
00050913
00078a63
01c42583
00048513
000780e7
06054c63
00c45783
0807f793
06079e63
03042583
00058c63
04040793
00f58663
00048513
ef5f50ef
02042823
04442583
00058863
00048513
ee1f50ef
04042223
d0df50ef
00041623
d09f50ef
00c12083
00812403
00412483
00090513
00012903
01010113
00008067
cd5f50ef
00c41783
f40786e3
f69ff06f
00c45783
fff00913
0807f793
f80786e3
01042583
00048513
e89f50ef
f7dff06f
040077b7
00050593
6747a503
ee5ff06f
fc010113
02c10313
02d12623
00030693
00112e23
02e12823
02f12a23
03012c23
03112e23
00612623
8f1fe0ef
01c12083
04010113
00008067
00050e13
04007537
fc010113
67452503
02810313
02c12423
02d12623
00058613
00030693
000e0593
00112e23
02e12823
02f12a23
03012c23
03112e23
00612623
8a1fe0ef
01c12083
04010113
00008067
fd010113
02812423
01312e23
01612823
02112623
02912223
03212023
01412c23
01512a23
00050b13
00058993
00060413
b00f90ef
00100793
02f51063
fff98793
0fe00713
00f76a63
0ff9f713
00e10623
00100913
02c0006f
05c40693
00098613
00c10593
000b0513
70c010ef
fff00793
00050913
0af50463
08050e63
00c14703
00000493
fff00a13
00a00a93
0280006f
00042783
00178693
00d42023
00e78023
00148493
00c10793
009787b3
0724f463
0007c703
00842783
fff78793
00f42423
fc07d8e3
01842683
00070593
00040613
000b0513
00d7c463
fb571ce3
854f50ef
fd4510e3
fff00913
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00090513
02012903
03010113
00008067
00098913
fd1ff06f
00c45783
0407e793
00f41623
fc1ff06f
00c61783
01279713
02074063
06462703
000026b7
00d7e7b3
000026b7
00d76733
00f61623
06e62223
eadff06f
fe010113
040077b7
00812c23
6747a403
00112e23
00058613
00050593
00040663
03842783
04078063
00c61783
01279713
02074063
06462703
000026b7
00d7e7b3
000026b7
00d76733
00f61623
06e62223
00040513
01812403
01c12083
02010113
e49ff06f
00a12423
00040513
00c12623
a45f50ef
00c12603
00812583
fadff06f
ff010113
00058713
00812423
00912223
00050413
040074b7
00060593
00070513
00112623
7804a823
5a5010ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
ff010113
00812423
00912223
00050413
040074b7
00058513
00112623
7804a823
5ad010ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
ff010113
00058713
00812423
00912223
00060593
00050413
040074b7
00068613
00070513
00112623
7804a823
5a5010ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
ff010113
00058713
00812423
00912223
00060593
00050413
040074b7
00068613
00070513
00112623
7804a823
fd9ed0ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
fe010113
01212823
0005a903
00812c23
00912a23
00112e23
01312623
01412423
00058413
00050493
04090263
00092983
02098863
0009aa03
000a0e63
000a2583
00058463
fbdff0ef
000a0593
00048513
a21f50ef
00098593
00048513
a15f50ef
00090593
00048513
a09f50ef
00040593
01812403
01c12083
01012903
00c12983
00812a03
00048513
01412483
02010113
9e1f506f
040077b7
6747a783
10a78a63
04c52583
fe010113
00912a23
00112e23
00812c23
01212823
01312623
00050493
04058063
00000913
08000993
012587b3
0007a403
00040e63
00040593
00042403
00048513
98df50ef
fe0418e3
04c4a583
00490913
fd391ce3
00048513
975f50ef
0404a583
00058663
00048513
965f50ef
1484a403
02040063
14c48913
01240c63
00040593
00042403
00048513
945f50ef
fe8918e3
0544a583
00058663
00048513
931f50ef
0384a783
04078663
03c4a783
00048513
000780e7
2e04a403
02040c63
00042583
00058663
00048513
e95ff0ef
00040593
01812403
01c12083
01012903
00c12983
00048513
01412483
02010113
8e1f506f
01c12083
01812403
01412483
01012903
00c12983
02010113
00008067
00008067
00862783
fd010113
01312e23
01412c23
02112623
02812423
02912223
03212023
01512a23
01612823
01712623
01812423
00062983
00060a13
14078863
0085a783
0005a703
00050a93
00058493
0d40006f
00c4d783
4807f693
08068a63
0144a603
0104a583
00161693
00c686b3
40b70433
01f6db13
00db0b33
00140713
401b5b13
01270733
000b0613
00eb7663
00070b13
00070613
4007f793
0a078a63
00060593
000a8513
854f90ef
00050c13
0a050e63
0104a583
00040613
935f90ef
00c4d783
b7f7f793
0807e793
00f49623
408b0733
008c0533
0164aa23
0184a823
00a4a023
00090b13
00e4a423
00090413
00040613
000b8593
a21f90ef
0084a783
0004a703
008a2683
416787b3
00870733
00f4a423
00e4a023
412686b3
00da2423
06068663
0049a903
0009ab83
00078b13
00898993
00078413
00070513
fe0904e3
f0f97ae3
00090b13
00090413
fa5ff06f
000a8513
d95fa0ef
00050c13
f6051ae3
0104a583
000a8513
f58f50ef
00c4d783
00c00713
00eaa023
0407e793
00f49623
000a2423
fff00513
0080006f
00000513
02c12083
02812403
000a2223
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
03010113
00008067
00c5d783
ed010113
11412c23
11612823
0fb12e23
12112623
12812423
12912223
13212023
11312e23
11512a23
11712623
11812423
11912223
11a12023
0807f793
00d12423
00058a13
00050b13
00060d93
00078663
0105a783
680784e3
00020737
04c10a93
00000813
57070713
00020c37
000204b7
000d8913
05512023
04012423
04012223
00012823
00012c23
00012e23
02012023
00012223
00e12623
6dcc0c13
6ec48493
00080993
000a8d93
00094703
1e070e63
00090413
02500693
2ad70863
00144703
00140413
fe071ae3
41240bb3
1d240e63
04412703
017989b3
012da023
00170713
017da223
05312423
04e12223
00700693
008d8d93
28e6c263
00412783
00044703
017787b3
00f12223
1a070063
00000693
00144603
00140913
02010da3
fff00e93
00012023
05a00b93
00900c93
02a00d13
00068413
00190913
fe060793
04fbe863
00c12703
00279793
00e787b3
0007a783
00078067
00012023
fd060793
00012683
00094603
00190913
00269713
00d70733
00171713
00e787b3
00f12023
fd060793
fcfcfee3
fe060793
fafbfce3
00040693
10060c63
08c10623
02010da3
00100b93
00100c93
08c10413
00000e93
0026ff93
000f8463
002b8b93
0846ff13
04412703
000f1863
00012783
41778d33
05a04ee3
03b14603
02060863
03b10613
00cda023
00170713
00100613
00198993
00cda223
05312423
04e12223
00700613
008d8d93
18e64c63
020f8863
03c10613
00cda023
00170713
00200613
00298993
00cda223
05312423
04e12223
00700613
008d8d93
12e64ee3
08000613
5acf0a63
419e8d33
6ba04c63
019989b3
00170713
008da023
019da223
05312423
04e12223
00700613
008d8793
76e64c63
0046f693
00068863
00012703
41770cb3
139048e3
00012403
01745463
000b8413
00412783
008787b3
00f12223
76099863
00094703
04012223
000a8d93
e00716e3
50099ce3
00ca5783
0407f793
580796e3
12c12083
12812403
00412503
12412483
12012903
11c12983
11812a03
11412a83
11012b03
10c12b83
10812c03
10412c83
10012d03
0fc12d83
13010113
00008067
000b0513
01d12a23
8adf80ef
00452783
00078513
02f12023
d79f10ef
00050793
000b0513
00f12e23
88df80ef
00852703
01c12783
01412e83
00e12c23
28079ee3
00094603
df9ff06f
00094603
02046413
dedff06f
00012703
00f12423
40e00733
00e12023
00094603
00446413
dd1ff06f
41240bb3
d72412e3
00044703
d95ff06f
04010613
000a0593
000b0513
ab9ff0ef
f20512e3
04812983
000a8d93
d65ff06f
04010613
000a0593
000b0513
03d12623
02d12423
03e12223
01f12a23
a89ff0ef
ee051ae3
04812983
04412703
02c12e83
02812683
02412f03
01412f83
000a8d93
e2dff06f
00812783
00040693
02010da3
0007a403
00478d13
3a0400e3
fff00713
00d12a23
2cee82e3
000e8613
00000593
00040513
01d12423
b50f90ef
00812e83
01412683
400506e3
40850cb3
01a12423
00000e93
0980006f
00812783
00040693
02010da3
0007a703
00478793
00f12423
08e10623
00100b93
00100c93
08c10413
d51ff06f
00040693
0206f713
1c070a63
00812783
00778793
ff87f793
0047a603
0007ac83
00878793
00f12423
00060b93
1e064263
fff00613
00068d13
00ce8863
017ce633
f7f6fd13
7a060a63
060b98e3
00900693
0796e4e3
030c8713
0ee107a3
000d0693
00100c93
0ef10413
000e8b93
019ed463
000c8b93
03b14703
00e03733
00eb8bb3
cd1ff06f
00812783
ffff86b7
8306c693
0007ac83
02d11e23
00478793
000216b7
00f12423
88c68793
00000b93
00246d13
00f12823
00200613
00000693
02d10da3
fff00693
16de8a63
017ce5b3
f7fd7693
4e059a63
260e9263
72061463
001d7c93
0f010413
f80c82e3
03000713
0ee107a3
0ef10413
f75ff06f
00812783
02047713
00478613
080716e3
01047713
200718e3
04047713
260712e3
20047693
200680e3
00812783
00c12423
0007a703
00412783
00f70023
b19ff06f
00094603
08046413
b99ff06f
00094603
06c00793
1af608e3
01046413
b85ff06f
00094603
06800793
1af606e3
04046413
b71ff06f
01046d13
020d7713
6a070a63
00812783
00100613
00778793
ff87f793
0007ac83
0047ab83
00878793
00f12423
f21ff06f
01046693
0206f713
6c070863
00812783
00778793
ff87f793
0007ac83
0047ab83
00878793
00f12423
bff6fd13
00000613
eedff06f
01046693
0206f713
e2071ae3
00812783
0106f613
0007a703
00478793
00f12423
62061463
0406f613
60060c63
01071c93
410cdc93
41fcdb93
000b8613
e20652e3
00068d13
02d00693
01903633
417008b3
02d10da3
fff00693
40c88bb3
41900cb3
00100613
e8de9ae3
00100693
e0d606e3
00200693
10d60463
0f010413
01db9793
007cf693
003cdc93
03068693
0197ecb3
003bdb93
fed40fa3
017ce7b3
00040593
fff40413
fc079ce3
001d7713
10070263
03000713
0ee68e63
ffe58593
0f010793
fee40fa3
40b78cb3
000d0693
00058413
dc9ff06f
00094603
00190713
15a602e3
fd060793
00070913
00000e93
a2fce0e3
00094603
002e9713
01d70eb3
001e9e93
00fe8eb3
fd060793
00190913
fefcf2e3
9fdff06f
02b00793
00094603
02f10da3
9e9ff06f
00812783
0007a703
00478793
00e12023
be0746e3
00094603
00f12423
9c9ff06f
00094603
00146413
9bdff06f
03b14783
00094603
9a0798e3
02000793
02f10da3
9a5ff06f
00100593
0ab600e3
00200593
00068d13
f0b610e3
01012683
0f010413
00fcf793
00f687b3
0007c703
004cdc93
01cb9793
0197ecb3
004bdb93
fee40fa3
017ce7b3
fff40413
fc079ce3
0f010793
40878cb3
000d0693
cddff06f
00012783
41778d33
a5a054e3
01000613
0ba65063
00812a23
00098793
000a0413
01000893
000d0a13
00700f13
00090d13
000e8993
00068913
00c0006f
ff0a0a13
0548da63
01078793
00170713
009da023
011da223
04f12423
04e12223
008d8d93
fcef5ee3
04010613
00040593
000b0513
de0ff0ef
3e051663
01000893
ff0a0a13
04812783
04412703
000a8d93
00700f13
fb48cae3
00090693
000d0913
000a0d13
00040a13
01412403
00098e93
00078993
01a989b3
00170713
009da023
01ada223
05312423
04e12223
00700613
008d8d93
98e650e3
04010613
000a0593
000b0513
03d12223
00d12a23
d68ff0ef
9c051ae3
02412e83
04812983
04412703
419e8d33
01412683
000a8d93
95a058e3
01000613
09a65863
00812a23
01000893
000a0413
00700e93
000d0a13
00090d13
00068913
00c0006f
ff0a0a13
0548da63
01098993
00170713
009da023
011da223
05312423
04e12223
008d8d93
fceedee3
04010613
00040593
000b0513
ce8ff0ef
2e051a63
01000893
ff0a0a13
04812983
04412703
000a8d93
00700e93
fb48cae3
00090693
000d0913
000a0d13
00040a13
01412403
01a989b3
00170713
009da023
01ada223
05312423
04e12223
00700613
008d8d93
88e65ce3
04010613
000a0593
000b0513
00d12a23
c7cff0ef
8e0514e3
04812983
04412703
01412683
000a8d93
86dff06f
04010613
000a0593
000b0513
00d12a23
c50ff0ef
8a051ee3
04812983
01412683
000a8793
869ff06f
04010613
000a0593
000b0513
c2cff0ef
88051ce3
04812983
87dff06f
00068d13
c71ff06f
01000613
0da65c63
000d0593
00090613
000d8793
000b8d13
000c8d93
00068b93
000a0913
00098693
01000893
00040993
00700293
01f12a23
03e12223
000e8c93
00060a13
00058413
00c0006f
ff040413
0488da63
01068693
00170713
0187a023
0117a223
04d12423
04e12223
00878793
fce2dee3
04010613
00090593
000b0513
b94ff0ef
4a051263
01000893
ff040413
04812683
04412703
000a8793
00700293
fa88cae3
01412f83
02412f03
00040613
000c8e93
000d8c93
00078d93
000a0793
00098413
00090a13
00068993
00078913
000b8693
000d0b93
00060d13
01a989b3
00170713
018da023
01ada223
05312423
04e12223
00700613
008d8d93
eae65663
04010613
000a0593
000b0513
03d12623
02d12423
03e12223
01f12a23
af8ff0ef
f6051263
04812983
04412703
02c12e83
02812683
02412f03
01412f83
000a8d93
e68ff06f
04010613
000a0593
000b0513
03d12423
02d12223
01e12a23
ab8ff0ef
f2051263
04812983
04412703
02812e83
02412683
01412f03
000a8d93
e90ff06f
01000693
04412703
0796d063
01000d13
00700413
00c0006f
ff0c8c93
059d5663
01098993
00170713
0187a023
01a7a223
05312423
04e12223
00878793
fce45ee3
04010613
000a0593
000b0513
a48ff0ef
ea051a63
ff0c8c93
04812983
04412703
000a8793
fb9d4ee3
019989b3
00170713
0187a023
0197a223
05312423
04e12223
00700793
e4e7d863
04010613
000a0593
000b0513
a00ff0ef
e6051663
04812983
e34ff06f
00040a13
e5cff06f
840e9ee3
000d0693
00000e93
00000c93
0f010413
85dff06f
2006f613
38061c63
41f75b93
00070c93
000b8613
809ff06f
00812783
010d7693
0007a703
00478793
00f12423
02069463
040d7693
00068c63
01071c93
010cdc93
00000b93
00100613
861ff06f
200d7693
32069e63
00070c93
00000b93
00100613
849ff06f
00812783
0106f613
0007a703
00478793
00f12423
02061263
0406f613
00060a63
01071c93
010cdc93
00000b93
925ff06f
2006f613
30061c63
00070c93
00000b93
911ff06f
400d7793
00000713
03312223
03412423
03212623
000c8993
000b8a13
01812903
0f010413
01d12a23
00078c93
00070b93
0240006f
00a00613
00000693
00098513
000a0593
511000ef
240a0c63
00050993
00058a13
00a00613
00000693
00098513
000a0593
2b0010ef
03050513
fea40fa3
001b8b93
fff40413
fa0c8ee3
00094683
fb769ae3
0ff00793
fafb86e3
140a1e63
00900793
1537ea63
0f010793
01212c23
01412e83
02412983
02812a03
02c12903
40878cb3
000d0693
ef8ff06f
01812783
00094603
b4078e63
0007c783
b4078a63
40046413
b4cff06f
0007a703
00412783
00c12423
41f7d693
00f72023
00d72223
aa4ff06f
00040d13
fc0ff06f
00021737
88c70793
00040693
00f12823
0206f713
06070263
00812783
00778793
ff87f793
0007ac83
0047ab83
00878793
00f12423
0016f593
00058e63
017ce5b3
00058a63
03000593
02b10e23
02c10ea3
0026e693
bff6fd13
00200613
ea8ff06f
00021737
8a070793
00040693
00f12823
0206f713
fa0712e3
00812783
0106f593
0007a703
00478793
00f12423
0a059463
0406f593
08058c63
01071c93
010cdc93
00000b93
f91ff06f
00040693
f40ff06f
00040513
9c4f10ef
01412683
00050c93
01a12423
00000e93
decff06f
04000593
854f80ef
00aa2023
00aa2823
18050263
04000793
00fa2a23
960ff06f
01c12783
02012583
00000b93
40f40433
00078613
00040513
8e5fa0ef
00194583
00a00613
00000693
00b03833
00098513
000a0593
01090933
335000ef
e29ff06f
2006f593
0a059663
00070c93
00000b93
ef9ff06f
00090a13
b58ff06f
00194603
02046413
00190913
9d0ff06f
00194603
20046413
00190913
9c0ff06f
00812783
0007a703
00412783
00c12423
00f72023
91cff06f
00600713
000e8c93
01d77463
00600c93
00021337
000c8b93
01a12423
8b430413
9f8ff06f
00900793
db37e4e3
df1ff06f
04010613
000a0593
000b0513
e71fe0ef
adcff06f
00812783
00c12423
0007a703
00412783
00f71023
8c0ff06f
0ff77c93
00000b93
e51ff06f
0ff77c93
00000b93
00100613
d10ff06f
01871c93
418cdc93
41fcdb93
000b8613
c70ff06f
0ff77c93
00000b93
dfcff06f
000e8c93
01a12423
00000e93
c90ff06f
00068d13
c74ff06f
fff00793
00f12223
a70ff06f
00812783
0007ae83
00478793
000ed463
fff00e93
00194603
00f12423
00070913
8c8ff06f
00c00793
00fb2023
fff00793
00f12223
a38ff06f
fe010113
00812c23
00912a23
040077b7
00112e23
1d87a783
00050413
00068493
02058263
000780e7
fff00793
02f50663
01c12083
01812403
01412483
02010113
00008067
00000613
00410593
000780e7
fff00793
fcf51ee3
0004a023
08a00793
01c12083
00f42023
01812403
01412483
02010113
00008067
fe010113
040077b7
00812c23
00912a23
00112e23
6747a483
040077b7
1d87a783
00060413
02050a63
00058613
00040693
00050593
00048513
000780e7
fff00793
02f50a63
01c12083
01812403
01412483
02010113
00008067
00060693
00410593
00000613
00048513
000780e7
fff00793
fcf51ae3
00042023
01c12083
01812403
08a00793
00f4a023
01412483
02010113
00008067
ff010113
00600513
00112623
368000ef
00100513
6e0000ef
000217b7
a2c7a703
14872783
04078c63
0047a703
01f00813
06e84e63
00271813
02050663
01078333
08c32423
1887a883
00100613
00e61633
00c8e8b3
1917a423
10d32423
00200693
02d50463
00170713
00e7a223
010787b3
00b7a423
00000513
00008067
14c70793
14f72423
fa5ff06f
18c7a683
00170713
00e7a223
00c6e6b3
18d7a623
010787b3
00b7a423
00000513
00008067
fff00513
00008067
2dc52783
00078663
00000513
00008067
ff010113
08000593
00812423
00112623
00050413
ccdf70ef
2ca42e23
02050463
08050793
00052023
00450513
fef51ce3
00000513
00c12083
00812403
01010113
00008067
fff00513
fedff06f
fe010113
00912a23
00112e23
00812c23
01f00793
00050493
02b7ea63
2dc52703
00058413
04070463
00241413
00870733
00072503
00c72023
01c12083
01812403
01412483
02010113
00008067
01c12083
01812403
01600793
00f52023
01412483
fff00513
02010113
00008067
08000593
00c12623
c21f70ef
2ca4ae23
00050713
02050063
00c12603
00050793
08050693
0007a023
00478793
fed79ce3
f8dff06f
fff00513
f95ff06f
ff010113
00912223
00112623
00812423
01f00793
00050493
0ab7ea63
2dc52783
00058413
04078463
00259713
00e787b3
0007a703
02070c63
00100693
06d70c63
fff00693
04d70863
00058513
0007a023
000700e7
00000513
00c12083
00812403
00412483
01010113
00008067
00048513
484000ef
00040613
00812403
00c12083
00050593
00048513
00412483
01010113
3fc0006f
00c12083
00812403
01600793
00f52023
00412483
00100513
01010113
00008067
00c12083
00812403
00412483
00000513
01010113
00008067
01600793
00f52023
fff00513
f81ff06f
01f00793
0cb7ea63
2dc52703
ff010113
00812423
00912223
00112623
00058413
00050493
06070063
00241793
00f70733
00072783
02078c63
fff00693
08d78663
00100693
06d78663
00040513
00072023
000780e7
00000513
00c12083
00812403
00412483
01010113
00008067
00c12083
00812403
00412483
00100513
01010113
00008067
08000593
a89f70ef
2ca4ae23
00050713
02050e63
00050793
08050693
0007a023
00478793
fed79ce3
f7dff06f
00c12083
00812403
00412483
00300513
01010113
00008067
00200513
f8dff06f
fff00513
f85ff06f
fff00513
00008067
ff010113
00912223
04007737
00112623
00812423
01f00793
67472483
0aa7e863
2dc4a783
00050413
04078263
00251713
00e787b3
0007a703
02070a63
00100693
06d70a63
fff00693
04d70663
0007a023
000700e7
00000513
00c12083
00812403
00412483
01010113
00008067
00048513
2c8000ef
00040613
00812403
00c12083
00050593
00048513
00412483
01010113
2400006f
00c12083
00812403
01600793
00f4a023
00100513
00412483
01010113
00008067
00c12083
00812403
00412483
00000513
01010113
00008067
01600793
00f4a023
fff00513
f81ff06f
ff010113
01212023
04007737
00112623
00812423
00912223
01f00793
67472903
02a7ee63
00050413
2dc92503
00058493
04050863
00241413
008507b3
0007a503
0097a023
00c12083
00812403
00412483
00012903
01010113
00008067
00c12083
00812403
01600793
00f92023
00412483
00012903
fff00513
01010113
00008067
08000593
00090513
8cdf70ef
2ca92e23
00050e63
00050793
08050713
0007a023
00478793
fee79ce3
f8dff06f
fff00513
f95ff06f
ff010113
040077b7
00812423
6747a403
00112623
2dc42783
00078c63
00000513
00c12083
00812403
01010113
00008067
08000593
00040513
869f70ef
2ca42e23
00050c63
08050793
00052023
00450513
fef51ce3
fc9ff06f
fff00513
fc5ff06f
ff010113
00912223
04007737
00112623
00812423
01f00793
67472483
0aa7ee63
2dc4a703
00050413
06070063
00241793
00f70733
00072783
02078c63
fff00693
08d78863
00100693
06d78863
00040513
00072023
000780e7
00000513
00c12083
00812403
00412483
01010113
00008067
00c12083
00812403
00412483
00100513
01010113
00008067
08000593
00048513
fb0f70ef
2ca4ae23
00050713
02050e63
00050793
08050693
0007a023
00478793
fed79ce3
f79ff06f
00c12083
00812403
00412483
00300513
01010113
00008067
00200513
f89ff06f
fff00513
f81ff06f
ff010113
00058713
00812423
00912223
00050413
040074b7
00060593
00070513
00112623
7804a823
160000ef
fff00793
00f50c63
00c12083
00812403
00412483
01010113
00008067
7904a783
fe0784e3
00c12083
00f42023
00812403
00412483
01010113
00008067
0d80006f
ff010113
00112623
00812423
03900893
00000073
00050413
00054c63
00c12083
00040513
00812403
01010113
00008067
40800433
ee9fd0ef
00852023
fff00413
fddff06f
05d00893
00000073
00054463
0000006f
ff010113
00812423
00050413
00112623
40800433
eb5fd0ef
00852023
0000006f
f7010113
08912223
08112623
00058493
08812423
05000893
00010593
00000073
00050413
02054463
00048513
00010593
0e0000ef
08c12083
00040513
08812403
08412483
09010113
00008067
40800433
e59fd0ef
00852023
fff00413
fcdff06f
00100513
00008067
f9010113
00810593
06112623
f8dff0ef
fff00793
00f50e63
00c12503
06c12083
00d55513
00157513
07010113
00008067
06c12083
00000513
07010113
00008067
ff010113
00112623
df9fd0ef
00c12083
01600793
00f52023
fff00513
01010113
00008067
ff010113
00112623
00812423
03e00893
00000073
00050413
00054c63
00c12083
00040513
00812403
01010113
00008067
40800433
da9fd0ef
00852023
fff00413
fddff06f
ff010113
0145a383
0185a283
01c5af83
0205af03
0305ae83
0405ae03
0385a303
0485a803
04c5a883
0585a603
00812623
00912423
0105a403
0085a483
01212223
0005a903
05c5a683
0685a703
06c5a783
01251023
00951123
00852223
00751423
00551523
01f51623
01e51723
01d52823
05c52623
04652423
01052c23
01152e23
02c52423
02d52623
00c12403
02e52c23
02f52e23
00812483
00412903
01010113
00008067
fd010113
01312e23
02112623
02812423
02912223
03212023
01412c23
01512a23
01612823
01712623
01812423
01912223
00050993
38069463
000207b7
00060a13
00050493
a1c78793
12c5f863
00010737
00058913
10e67863
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
02000693
00e787b3
40f68733
00f68c63
00e59933
00f9d7b3
00e61a33
0127e933
00e994b3
010a5a93
000a8593
00090513
010a1b13
fadef0ef
010b5b13
00050593
00050993
000b0513
f6def0ef
00050413
000a8593
00090513
fd1ef0ef
01051513
0104d713
00a76733
00098913
00877e63
01470733
fff98913
01476863
00877663
ffe98913
01470733
40870433
000a8593
00040513
f4def0ef
00050593
00050993
000b0513
f11ef0ef
00050b13
000a8593
00040513
f75ef0ef
01049713
01051513
01075713
00a76733
00098693
01677c63
00ea0733
fff98693
01476663
01677463
ffe98693
01091793
00d7e7b3
00000913
1200006f
010006b7
01000713
eed66ce3
01800713
ef1ff06f
00061463
00100073
00010737
12e67c63
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
02000693
00e787b3
40f68733
12f69263
40c589b3
00100913
010a5b13
000b0593
00098513
010a1b93
e89ef0ef
010bdb93
00050593
00050c13
000b8513
e49ef0ef
00050a93
000b0593
00098513
eadef0ef
01051513
0104d713
00a76733
000c0993
01577e63
01470733
fffc0993
01476863
01577663
ffec0993
01470733
41570433
000b0593
00040513
e29ef0ef
00050593
00050a93
000b8513
dedef0ef
00050b93
000b0593
00040513
e51ef0ef
01049713
01051513
01075713
00a76733
000a8693
01777c63
00ea0733
fffa8693
01476663
01777463
ffea8693
01099793
00d7e7b3
02c12083
02812403
02412483
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00090593
00078513
02012903
03010113
00008067
010006b7
01000713
ecd668e3
01800713
ec9ff06f
00e61a33
00f5d933
010a5b93
00e595b3
00f9d7b3
00b7eab3
00e994b3
000b8593
00090513
010a1993
d59ef0ef
0109d993
00050593
00050b13
00098513
d19ef0ef
00050413
000b8593
00090513
d7def0ef
01051513
010ad713
00a76733
000b0913
00877e63
01470733
fffb0913
01476863
00877663
ffeb0913
01470733
40870433
000b8593
00040513
cf9ef0ef
00050593
00050b13
00098513
cbdef0ef
00050993
000b8593
00040513
d21ef0ef
010a9793
01051513
0107d793
00a7e7b3
000b0713
0137fe63
014787b3
fffb0713
0147e863
0137f663
ffeb0713
014787b3
01091913
413789b3
00e96933
e01ff06f
1ed5ec63
000107b7
04f6f463
1006b513
00154513
00351513
000207b7
00a6d733
a1c78793
00e787b3
0007c703
02000793
00a70733
40e78933
02e79663
00100793
e8b6e2e3
00c9b7b3
0017c793
e79ff06f
010007b7
01000513
fcf6e0e3
01800513
fb9ff06f
012696b3
00e65b33
00db6b33
00e5da33
010b5c13
00e9d733
012595b3
00b76ab3
000a0513
000c0593
010b1b93
012614b3
010bdb93
bfdef0ef
00050593
00050c93
000b8513
bc1ef0ef
00050413
000c0593
000a0513
c25ef0ef
01051513
010ad693
00a6e6b3
000c8a13
0086fe63
016686b3
fffc8a13
0166e863
0086f663
ffec8a13
016686b3
40868433
000c0593
00040513
ba1ef0ef
00050593
00050c93
000b8513
b65ef0ef
00050b93
000c0593
00040513
bc9ef0ef
010a9713
01051513
01075713
00a76733
000c8693
01777e63
01670733
fffc8693
01676863
01777663
ffec8693
01670733
010a1793
00010e37
00d7e7b3
fffe0313
41770833
0067f733
0064f333
0107de93
0104d493
00070513
00030593
af5ef0ef
00050893
00048593
00070513
ae5ef0ef
00050713
00030593
000e8513
ad5ef0ef
00050313
00048593
000e8513
ac5ef0ef
00670733
0108d693
00d70733
00677463
01c50533
01075693
00a686b3
02d86663
bcd81ce3
00010637
fff60613
00c77733
01071713
00c8f8b3
012996b3
01170733
00000913
cce6fce3
fff78793
badff06f
00000913
00000793
cc5ff06f
fd010113
02812423
02912223
02112623
03212023
01312e23
01412c23
01512a23
01612823
01712623
01812423
01912223
01a12023
00050413
00058493
24069c63
000207b7
00060a13
a1c78793
12c5fe63
00010737
12e67063
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
00e787b3
02000713
40f70933
00f70c63
012595b3
00f557b3
01261a33
00b7e4b3
01251433
010a5a93
000a8593
010a1b13
00048513
9edef0ef
010b5b13
000b0593
9b5ef0ef
00050993
000a8593
00048513
a19ef0ef
01051513
01045793
00a7e7b3
0137fa63
014787b3
0147e663
0137f463
014787b3
413784b3
000a8593
00048513
9a1ef0ef
000b0593
96def0ef
00050993
000a8593
00048513
9d1ef0ef
01041413
01051513
01045413
00a46433
01347a63
01440433
01446663
01347463
01440433
41340433
01245533
00000593
02c12083
02812403
02412483
02012903
01c12983
01812a03
01412a83
01012b03
00c12b83
00812c03
00412c83
00012d03
03010113
00008067
010006b7
01000713
eed664e3
01800713
ee1ff06f
00061463
00100073
00010737
0ee67663
10063713
00174713
00371713
00e656b3
00d787b3
0007c783
40c584b3
00e787b3
02000713
40f70933
ecf70ae3
01261a33
00f5dbb3
010a5b13
00f557b3
012595b3
00b7e9b3
01251433
000b0593
010a1a93
000b8513
8a5ef0ef
010ada93
000a8593
86def0ef
00050493
000b0593
000b8513
8d1ef0ef
01051513
0109d713
00a76733
00977a63
01470733
01476663
00977463
01470733
409704b3
000b0593
00048513
859ef0ef
000a8593
825ef0ef
00050a93
000b0593
00048513
889ef0ef
01099793
01051513
0107d793
00a7e7b3
0157fa63
014787b3
0147e663
0157f463
014787b3
415784b3
e19ff06f
010006b7
01000713
f0d66ee3
01800713
f15ff06f
ead5e4e3
000107b7
04f6fe63
1006b793
0017c793
00379793
00020737
00f6d833
a1c70713
01070733
00074983
00f989b3
02000793
41378933
05379063
00b6e463
00c56c63
40c50633
40d586b3
00c535b3
40b684b3
00060413
00040513
00048593
e49ff06f
01000737
01000793
fae6e6e3
01800793
fa5ff06f
012696b3
01365b33
00db6b33
0135d4b3
01355a33
012595b3
010b5c93
00ba6a33
01251ab3
000c8593
00048513
010b1c13
01261bb3
010c5c13
f4cef0ef
00050593
00050d13
000c0513
f10ef0ef
00050413
000c8593
00048513
f74ef0ef
01051513
010a5793
00a7e7b3
000d0493
0087fe63
016787b3
fffd0493
0167e863
0087f663
ffed0493
016787b3
40878433
000c8593
00040513
ef0ef0ef
00050593
00050d13
000c0513
eb4ef0ef
000c8593
00050c13
00040513
f18ef0ef
010a1593
01051513
0105d593
00a5e5b3
000d0793
0185fe63
016585b3
fffd0793
0165e863
0185f663
ffed0793
016585b3
00010eb7
01049493
00f4e4b3
fffe8793
00f4f8b3
00fbf7b3
41858733
0104d493
010bde13
00088513
00078593
e44ef0ef
00050813
000e0593
00088513
e34ef0ef
00050893
00078593
00048513
e24ef0ef
00050313
000e0593
00048513
e14ef0ef
01085793
006888b3
011787b3
00050613
0067f463
01d50633
0107d693
00c686b3
00010637
fff60613
00c7f7b3
01079793
00c87833
010787b3
00d76663
00d71e63
00fafc63
41778633
00c7b7b3
016787b3
40f686b3
00060793
40fa87b3
00fabab3
40d705b3
415585b3
013599b3
0127d7b3
00f9e533
0125d5b3
c71ff06f
00c52783
0005af03
0045af83
0085a283
00c5a583
00008737
0107d693
fff70713
01079813
01059e93
01f7d613
00e6f6b3
0105d793
00052883
00452303
00852e03
ff010113
01085813
010ede93
00e7f7b3
01f5d593
02e69063
0068e733
01c76733
01076733
00100513
04071a63
04d79863
0080006f
00e79c63
01ff6733
00576733
01d76733
00100513
02071a63
00100513
02d79663
03e89463
03f31263
025e1063
01d81e63
02b60063
00079a63
0068e533
01c56533
01056533
00a03533
01010113
00008067
00000513
ff5ff06f
00052f83
00452803
00852e03
00c52503
00c5a683
000087b7
01055613
fff78793
01069313
0106d713
0005a283
0045a883
0085ae83
00f67633
01051593
ff010113
0105d593
01f55513
01035313
00f77733
01f6d693
00f61e63
01f867b3
01c7e7b3
00b7e7b3
0c078863
ffe00513
0640006f
00f71a63
0112e7b3
01d7e7b3
0067e7b3
fe0794e3
0a061a63
01f867b3
01c7e7b3
00b7e7b3
0017b793
00071a63
0112ef33
01df6f33
006f6f33
060f0a63
00079c63
00a69463
02c75263
04050e63
fff00513
0100006f
fff00513
00068463
00068513
01010113
00008067
00e65663
fe051ae3
fddff06f
fcb36ae3
02659e63
fdcee6e3
03de1e63
fd08e2e3
01181463
fbf2eee3
fd186ee3
01181463
fc5feae3
00000513
fc1ff06f
00100513
fb9ff06f
fe0798e3
f99ff06f
fa65ece3
fe5ff06f
fbde68e3
fddff06f
f4c700e3
f6071ce3
00000793
f5dff06f
00052f83
00452803
00852e03
00c52503
00c5a683
000087b7
01055613
fff78793
01069313
0106d713
0005a283
0045a883
0085ae83
00f67633
01051593
ff010113
0105d593
01f55513
01035313
00f77733
01f6d693
00f61e63
01f867b3
01c7e7b3
00b7e7b3
0c078863
00200513
0640006f
00f71a63
0112e7b3
01d7e7b3
0067e7b3
fe0794e3
0a061a63
01f867b3
01c7e7b3
00b7e7b3
0017b793
00071a63
0112ef33
01df6f33
006f6f33
060f0a63
00079c63
00a69463
02c75263
04050e63
fff00513
0100006f
fff00513
00068463
00068513
01010113
00008067
00e65663
fe051ae3
fddff06f
fcb36ae3
02659e63
fdcee6e3
03de1e63
fd08e2e3
01181463
fbf2eee3
fd186ee3
01181463
fc5feae3
00000513
fc1ff06f
00100513
fb9ff06f
fe0798e3
f99ff06f
fa65ece3
fe5ff06f
fbde68e3
fddff06f
f4c700e3
f6071ce3
00000793
f5dff06f
f6010113
09312623
00c5a983
0005a783
0085a683
08912a23
00050493
0045a503
01099713
09412423
09512223
00c62a03
00062a83
09612023
07712e23
00862b03
00462b83
00008637
09212823
01075713
0109d913
fff60613
05312623
08112e23
08812c23
07812c23
07912a23
07a12823
07b12623
04f12023
04a12223
04d12423
00f12823
00a12a23
00d12c23
00e12e23
00c97933
01f9d993
580906e3
6ac902e3
000107b7
00f76733
00e12e23
01010613
01c10793
0007a703
ffc7a683
ffc78793
00371713
01d6d693
00d76733
00e7a223
fef612e3
01012783
00379793
00f12823
ffffc7b7
00178793
00f90933
00000c13
010a1513
00008737
010a5793
01055513
fff70713
05412623
05512023
05712223
05612423
03512023
03712223
03612423
02a12623
00e7f7b3
01fa5a13
62078ee3
00e79463
7510006f
00010737
00e56533
02a12623
02010593
02c10713
00072683
ffc72603
ffc70713
00369693
01d65613
00c6e6b3
00d72223
fee592e3
02012703
00371713
02e12023
ffffc737
00170713
00e787b3
00000693
012787b3
00f12423
00178c93
002c1793
00d7e7b3
00a00713
0149c433
00f75463
74d0006f
00200713
00f75463
6fd0006f
fff78793
00100713
00f76463
7950006f
01012283
02012f83
00010337
fff30793
00f2f833
00fff7b3
0102de93
010fd713
00080513
00078593
850ef0ef
00050e13
00070593
00080513
840ef0ef
00050813
00078593
000e8513
830ef0ef
00050893
00070593
000e8513
820ef0ef
010e5713
01180833
01070733
00050793
01177463
006507b3
01075693
00f687b3
00010337
02412e83
04f12223
fff30793
00f77733
01071713
00fe7533
00a70533
00fef833
00f2f733
04a12023
0102d893
010edf13
00070513
00080593
fc1ee0ef
00050e13
000f0593
00070513
fb1ee0ef
00050713
00080593
00088513
fa1ee0ef
00050813
000f0593
00088513
f91ee0ef
010e5893
01070733
00e888b3
00050a13
0108f463
00650a33
01412f03
0108d713
00f8f8b3
00fe7533
00e12623
01089893
00ff7733
00fff7b3
00a888b3
010f5393
010fd313
00070513
00078593
f41ee0ef
00050813
00030593
00070513
f31ee0ef
00050713
00078593
00038513
f21ee0ef
00050e13
00030593
00038513
f11ee0ef
01085313
01c70733
00e30333
00050793
01c37663
00010737
00e507b3
00010e37
fffe0593
01035b93
00b37333
00b87833
00bf7933
00bef3b3
01031313
00fb8bb3
01030333
010ed793
010f5813
00090513
00038593
eb9ee0ef
00050713
00078593
00090513
ea9ee0ef
00050913
00038593
00080513
e99ee0ef
00050393
00078593
00080513
e89ee0ef
01075813
007906b3
00d80833
00050793
00787463
01c507b3
00010e37
fffe0593
02812383
01085b13
00b87833
00b77733
01081813
00b2f933
00e80833
00b3f733
00fb0b33
0102dc13
0103da93
00090513
00070593
e31ee0ef
00050793
000a8593
00090513
e21ee0ef
00050993
00070593
000c0513
e11ee0ef
00050913
000a8593
000c0513
e01ee0ef
0107d713
012986b3
00d70733
01277463
01c50533
00010d37
fffd0913
01812e03
01075a93
01277733
0127f7b3
01071713
00f70733
012e77b3
012ff933
00aa8ab3
010e5d93
010fdc13
00078513
00090593
dadee0ef
00050993
000c0593
00078513
d9dee0ef
00050793
00090593
000d8513
d8dee0ef
00050913
000c0593
000d8513
d7dee0ef
012787b3
0109d693
00d787b3
0127f463
01a50533
00010937
fff90593
04412603
0107d693
00b7f7b3
01079793
00b9f9b3
013789b3
00c12783
00c88633
011638b3
011787b3
00660633
01478a33
017a07b3
04c12223
00663633
00c78333
00a68533
0177b7b3
010306b3
00c33333
011a3a33
0067e7b3
014787b3
0106b833
016787b3
01078a33
00e686b3
00e6b733
015a08b3
00e88333
013686b3
00a30633
04d12423
0136b6b3
00d609b3
010a3a33
0167b7b3
0158b8b3
00e33333
02c12803
05312623
0147e7b3
00d9b9b3
0068e8b3
00a63633
01366633
011787b3
00c787b3
04f12823
0102da13
00b877b3
00b2f2b3
01085993
00028513
00078593
c81ee0ef
00050713
00098593
00028513
c71ee0ef
00050893
00078593
000a0513
c61ee0ef
00050313
00098593
000a0513
c51ee0ef
01075613
006888b3
01160633
00050793
00667463
012507b3
01065a13
000102b7
01c12883
00fa0a33
fff28793
00f67633
00f77733
01061613
00e60333
00f8f933
010fd713
00ffffb3
0108d993
00090513
000f8593
bf9ee0ef
00050793
00070593
00090513
be9ee0ef
00050913
000f8593
00098513
bd9ee0ef
00050f93
00070593
00098513
bc9ee0ef
0107d693
01f90933
012686b3
00050713
01f6f463
00550733
00010fb7
ffff8613
0106d993
00c6f6b3
01069693
00c7f7b3
00cf7933
00c3f2b3
00e989b3
00f68b33
010f5713
0103da93
00090513
00028593
b75ee0ef
00050793
000a8593
00090513
b65ee0ef
00050913
00028593
00070513
b55ee0ef
00050293
000a8593
00070513
b45ee0ef
0107d713
005906b3
00d70733
00577463
01f50533
000102b7
fff28693
01075913
00d77733
00d7f7b3
00de7ab3
00deffb3
01071713
00a90933
00f70733
010e5d13
010edc13
000a8513
000f8593
af5ee0ef
00050793
000c0593
000a8513
ae5ee0ef
00050b93
000f8593
000d0513
ad5ee0ef
00050a93
000c0593
000d0513
ac5ee0ef
0107df93
015b86b3
00df8fb3
015ff463
00550533
00010ab7
fffa8293
010fdb93
005fffb3
0057f7b3
010f9f93
00ff8fb3
04c12783
00ab8bb3
00f307b3
0067b633
05012303
016787b3
0167b6b3
006a0333
00c30d33
013d0b33
00db0c33
00e787b3
00e7b733
012c05b3
00e58533
01f787b3
04f12623
01433333
01f7b7b3
00cd3d33
01750fb3
013b3b33
00dc3c33
00ff8db3
00e53533
01a36333
018b6b33
0125b5b3
00a5e5b3
05b12823
01630333
00fdbdb3
017fbfb3
00b30333
01bfefb3
01f307b3
005e7333
0053f2b3
04f12a23
010e5913
0103d713
00030513
00028593
9e5ee0ef
00050793
00070593
00030513
9d5ee0ef
00050313
00028593
00090513
9c5ee0ef
00050f93
00070593
00090513
9b5ee0ef
0107d613
01f30333
00660633
00050713
01f67463
01550733
01065993
00010fb7
00e989b3
ffff8713
00e67633
01061613
00e7f7b3
010f5a13
00ef7f33
00e87733
00f607b3
01085913
000f0513
00070593
961ee0ef
00050313
00090593
000f0513
951ee0ef
00050f13
00070593
000a0513
941ee0ef
00050293
00090593
000a0513
931ee0ef
01035693
005f0f33
01e686b3
00050713
0056f463
01f50733
000102b7
fff28613
0106d913
00c6f6b3
00c37333
01069693
00668a33
010edf13
00c8f333
00cefeb3
00e90933
00030513
0108d713
000e8593
8ddee0ef
00050f93
000f0593
00030513
8cdee0ef
00050a93
000e8593
00070513
8bdee0ef
00050313
000f0593
00070513
8adee0ef
00050713
010fdf13
006a8533
00af0f33
006f7463
00570733
010f5293
00010337
00e282b3
fff30713
00ef7f33
00efffb3
010f1f13
01ff0f33
010e5a93
00e87fb3
00ee7e33
01085b13
000e0513
000f8593
859ee0ef
00050e93
000b0593
000e0513
849ee0ef
00050713
000f8593
000a8513
839ee0ef
00050f93
000b0593
000a8513
829ee0ef
01f70733
010ed693
00d70733
01f77463
00650533
00010337
fff30593
01075f93
00b77733
00befeb3
00b8fb33
0103db93
01071713
00b3f3b3
00af8fb3
01d70733
0108de13
000b0513
00038593
fd8ee0ef
00050a93
000b8593
000b0513
fc8ee0ef
00050b13
00038593
000e0513
fb8ee0ef
00050393
000b8593
000e0513
fa8ee0ef
010ade93
007b06b3
00de8eb3
007ef463
00650533
05012583
00010e37
fffe0313
00b785b3
00f5b633
05412783
014585b3
0145b6b3
00f987b3
00c78bb3
012b8a33
00da0b33
01e585b3
010ed393
006efeb3
00a383b3
006afab3
005b0533
04b12823
010e9e93
01e5b5b3
015e8eb3
00cbbbb3
00b50ab3
00db3b33
0137b7b3
012a3a33
00ea8f33
0177e7b3
00babab3
016a6a33
00553533
01556533
014787b3
00a787b3
00ef3733
01f787b3
00e785b3
01df0f33
007586b3
05e12a23
01df3f33
01e68633
00e5b5b3
04c12c23
01f7b7b3
01e63633
0076b6b3
00b7e7b3
00c6e6b3
00d787b3
04f12e23
0108df13
01085793
0068f8b3
00687833
00088513
00080593
ea8ee0ef
00050e93
00078593
00088513
e98ee0ef
00050713
00080593
000f0513
e88ee0ef
00050813
00078593
000f0513
e78ee0ef
010ed793
01070733
00e787b3
00050693
0107f463
01c506b3
05812603
0067f733
05c12583
01071713
006efeb3
01d70733
00c70633
0107d793
00b787b3
00e63733
00e787b3
00d78533
04412703
04012783
04a12e23
04c12c23
00f76733
04812783
05010593
00f76733
04c12783
00d79793
00e7e7b3
04010713
00c72683
01072603
00470713
0136d693
00d61613
00c6e6b3
fed72e23
fee592e3
04812683
04012703
00f037b3
02d12c23
04412683
00e7e7b3
04c12703
02d12a23
001006b7
02e12e23
02f12823
00d77733
4e070463
01f79793
03010713
03c10593
00072683
00472603
00470713
0016d693
01f61613
00c6e6b3
fed72e23
fee592e3
03c12703
00f037b3
00175713
02e12e23
03012703
00f767b3
02f12823
000047b7
fff78793
00fc87b3
4af05863
03012703
00777693
04068463
00f77693
00400613
02c68e63
03412683
00470713
02e12823
00473713
00d706b3
02d12a23
00e6b6b3
03812703
00e68733
02e12c23
00d73733
03c12683
00d70733
02e12e23
03c12703
001006b7
00d776b3
00068e63
fff007b7
fff78793
00f77733
000047b7
02e12e23
00fc87b3
03010713
03c10593
00072683
00472603
00470713
0036d693
01d61613
00c6e6b3
fed72e23
feb712e3
000086b7
ffe68613
03c12703
3ef64463
00375713
02e12e23
01179793
0117d793
00f41413
00f46433
03012783
03c12703
04811723
00f4a023
03412783
04e11623
09c12083
00f4a223
03812783
09812403
09012903
00f4a423
04c12783
08c12983
08812a03
00f4a623
08412a83
08012b03
07c12b83
07812c03
07412c83
07012d03
06c12d83
00048513
09412483
0a010113
00008067
00a7e633
00d66633
00e66633
12060663
08070463
00070513
d4cee0ef
00050413
ff440593
4055d793
01f5f593
40f00733
08058e63
00271713
00c70693
02000513
01010893
40b50533
00d886b3
40e00733
0ad89463
fff78613
00279793
01010713
05078793
00e787b3
01012703
00b71733
fae7a823
00160613
ffffc937
00261613
00000593
01010513
01190913
de4ee0ef
40890933
a34ff06f
00068a63
00068513
cc4ee0ef
02050413
f79ff06f
00050863
cb4ee0ef
04050413
f69ff06f
00078513
ca4ee0ef
06050413
f59ff06f
01c10693
00271713
00300613
00e685b3
0005a583
fff60613
ffc68693
00b6a223
fef656e3
fff78613
f81ff06f
0006a603
ffc6a803
00e68333
00b61633
00a85833
01066633
00c32023
ffc68693
f39ff06f
00a7e7b3
00d7e7b3
00e7e7b3
00300c13
9a079063
00200c13
998ff06f
00000913
00100c13
98cff06f
017ae7b3
0167e7b3
00a7e7b3
12078863
08050263
c0cee0ef
00050413
ff440593
4055d793
01f5f593
40f00733
0a058063
00271713
00c70693
02000513
02010893
40b50533
00d886b3
40e00733
0ad89663
fff78613
00279793
01010713
05078793
00e787b3
02012703
00b71733
fce7a023
00160613
00261613
00000593
02010513
cacee0ef
ffffc7b7
01178793
408787b3
98cff06f
000b0a63
000b0513
b84ee0ef
02050413
f79ff06f
000b8a63
000b8513
b70ee0ef
04050413
f65ff06f
000a8513
b60ee0ef
06050413
f55ff06f
02c10693
00271713
00300613
00e685b3
0005a583
fff60613
ffc68693
00b6a223
fef656e3
fff78613
f7dff06f
0006a603
ffc6a803
00e68333
00b61633
00a85833
01066633
00c32023
ffc68693
f35ff06f
017aeab3
016aeab3
00aaeab3
00300693
000a8463
8f0ff06f
00200693
8e8ff06f
00000793
00100693
8dcff06f
00100713
00f717b3
5307f713
04071663
0887f713
08071863
2407f793
00079463
8f8ff06f
000087b7
02f12e23
02012c23
02012a23
02012823
fff78793
00000413
cb9ff06f
00f00713
fce78ee3
00b00713
04e78a63
00098413
01012783
02f12823
01412783
02f12a23
01812783
02f12c23
01c12783
02f12e23
00200793
26fc0e63
00300793
fafc00e3
00100793
bafc12e3
02012e23
02012c23
02012a23
02012823
2180006f
000a0413
02012783
00068c13
02f12823
02412783
02f12a23
02812783
02f12c23
02c12783
fadff06f
00812c83
b61ff06f
02012e23
02012c23
02012a23
02012823
fff68793
c11ff06f
00100713
40f707b3
07400713
1cf74463
03010993
4057d513
00098693
00000913
00000713
04a71263
01f7f793
00251693
04079663
00300613
00098793
00000713
40a60633
00d785b3
0005a583
00170713
00478793
feb7ae23
fee656e3
00400793
40a78533
0780006f
0006a603
00170713
00468693
00c96933
fadff06f
05068713
01010613
00c70733
fd072703
02000593
40f585b3
00b71733
00e96933
00300713
00d986b3
00098893
00000813
40a70733
00468693
0ce84263
00400693
00271713
40a68533
05070713
01010693
00d70733
03c12683
00f6d7b3
fcf72823
00400a13
40aa0633
00251513
00261613
00000593
00a98533
a04ee0ef
03012703
012037b3
00e7e7b3
02f12823
0077f713
04070263
00f7f713
03470e63
03412703
00478793
02f12823
0047b793
00e78733
02e12a23
00f73733
03812783
00f707b3
02f12c23
00e7b7b3
03c12703
00e787b3
02f12e23
03c12703
000807b7
00e7f7b3
04078063
02012e23
02012c23
02012a23
02012823
00100793
a99ff06f
ffc6a603
0006a303
00180813
00f65633
00b31333
00666633
00c8a023
00488893
f19ff06f
00c98693
0009a783
0049a703
00498993
0037d793
01d71713
00e7e7b3
fef9ae23
fed992e3
03c12783
0037d793
02f12e23
00000793
a3dff06f
03412783
03012703
00f76733
03812783
00f76733
03c12783
00f76733
00000793
a0070ce3
02012e23
02012c23
02012a23
02012823
a05ff06f
000087b7
02012e23
02012c23
02012a23
02012823
fff78793
9e9ff06f
f9010113
0085a783
05312e23
00c5a983
0005a683
0045a703
05412c23
05712623
00050a13
02f12c23
00f12c23
00062883
01099793
00462503
00862583
00c62b83
06812423
0107d793
00199413
02d12823
03312e23
00d12823
06112623
06912223
07212023
05512a23
05612823
05812423
05912223
02e12a23
00e12a23
00f12e23
01145413
01f9d993
01010813
01c10693
0006a783
ffc6a703
ffc68693
00379793
01d75713
00e7e7b3
00f6a223
fed812e3
01012903
010b9793
001b9b13
00391913
0107d793
02a12a23
03712e23
02a12223
01212823
03112823
02b12c23
03112023
02b12423
02f12623
011b5b13
01fbdb93
02010513
02c10713
00072783
ffc72603
ffc70713
00379793
01d65613
00c7e7b3
00f72223
fee512e3
02012483
000087b7
fff78793
00349493
02912023
02fb1063
02812603
02412783
00c7e7b3
02c12603
00c7e7b3
0097e7b3
00079463
001bcb93
416405b3
113b94e3
2eb05463
01412c03
01812b83
01c12a83
0a0b1a63
02412603
02812783
02c12803
00f666b3
0106e6b3
0096e6b3
00069e63
03212823
03812a23
03712c23
03512e23
00058413
2ec0006f
fff58693
04069863
009904b3
01860633
02912823
0124b4b3
00960733
02e12a23
01863633
00973733
00e66633
017787b3
00c78733
02e12c23
0177b7b3
00c73733
00e7e7b3
01580833
010787b3
00100413
19c0006f
000087b7
fff78793
f8f586e3
07400793
04d7da63
02012623
02012423
02012223
00100793
11c0006f
000087b7
fff78793
00f41c63
03212823
03812a23
03712c23
03512e23
2500006f
02c12783
000806b7
00d7e7b3
02f12623
07400793
fab7cce3
00058693
4056d793
00070593
00000493
00000613
02f61e63
01f6f693
00279593
04069263
00300613
40f60633
00b70833
00082803
00168693
00470713
ff072e23
fed656e3
00400713
40f707b3
06c0006f
0005a803
00160613
00458593
0104e4b3
fb5ff06f
04058613
00260633
fe062603
02000893
40d888b3
01161633
00c4e4b3
00300613
00b505b3
00000313
40f60633
00458593
12c34a63
00400713
00261613
40f707b3
04060713
00270633
02c12703
00d75733
fee62023
00400613
40f60633
00279793
00f50533
00261613
00000593
daded0ef
02012703
009037b3
00f767b3
02f12023
02012783
02412703
00f907b3
00ec0733
02f12823
0127b7b3
00f706b3
02d12a23
00f6b6b3
02812783
01873733
00d76733
00fb87b3
00e786b3
02d12c23
00e6b6b3
02c12703
0177b7b3
00d7e7b3
00ea8733
00e787b3
00080737
02f12e23
00e7f733
0e070863
fff80737
fff70713
00e7f7b3
02f12e23
03012783
00140413
03c10593
01f79713
03010793
0007a683
0047a603
00478793
0016d693
01f61613
00c6e6b3
fed7ae23
feb792e3
03c12783
0017d793
02f12e23
00e037b3
03012703
00f767b3
02f12823
000087b7
fff78793
08f41263
02012e23
02012c23
02012a23
02012823
0700006f
ffc5a803
0005ae03
00130313
00d85833
011e1e33
01c86833
01072023
00470713
ea9ff06f
02412a83
02812b83
02c12c03
40058063
408b0633
20041a63
01412703
01812783
01c12503
00f765b3
00a5e5b3
0125e5b3
18059063
02912823
03512a23
03712c23
03812e23
00060413
03012783
0077f713
04070463
00f7f713
00400693
02d70e63
03412703
00478793
02f12823
0047b793
00e78733
02e12a23
00f73733
03812783
00f707b3
02f12c23
00e7b7b3
03c12703
00e787b3
02f12e23
03c12783
00080737
00e7f733
02070463
00008737
00140413
fff70713
00e41463
0100106f
fff80737
fff70713
00e7f7b3
02f12e23
03010793
03c10613
0007a703
0047a683
00478793
00375713
01d69693
00d76733
fee7ae23
fef612e3
03c12703
000086b7
fff68793
00375713
02e12e23
02f41a63
03412603
03012783
00c7e7b3
03812603
00c7e7b3
00e7e7b3
00078c63
02d12e23
02012c23
02012a23
02012823
00000993
03c12783
01141413
01145413
00f11623
03012783
00f99993
0089e9b3
00fa2023
03412783
01311723
06c12083
00fa2223
03812783
06812403
06412483
00fa2423
00c12783
06012903
05c12983
00fa2623
05412a83
05012b03
04c12b83
04812c03
04412c83
000a0513
05812a03
07010113
00008067
fff60893
04089663
00990933
01570733
03212823
00993933
012706b3
02d12a23
01573733
0126b6b3
00d76733
017787b3
00e786b3
02d12c23
0177b7b3
00e6b6b3
00d7e7b3
01850533
00a787b3
bb1ff06f
000087b7
fff78793
e2f606e3
07400793
0517dc63
00012e23
00012c23
00012a23
00100793
1640006f
000087b7
fff78793
00fb1e63
02912823
03512a23
03712c23
03812e23
000b0413
e01ff06f
01c12783
00080737
00e7e7b3
00f12e23
07400793
fac7cae3
00060893
41f8d793
01f7f793
011787b3
4057d793
00068613
00000413
00000713
04f74663
00078593
0007d463
00000593
01f8f513
00279613
04051463
00300593
00000713
40f585b3
00c68533
00052503
00170713
00468693
fea6ae23
fee5d6e3
00400713
40f707b3
08c0006f
00062583
00170713
00460613
00b46433
fa5ff06f
80000737
01f70713
00e8f733
00075863
fff70713
fe076713
00170713
00259593
02000893
40e888b3
04058713
002705b3
fd05a703
00c80633
00000313
01171733
00e46433
00300713
40f70733
00460613
0ae34a63
00400693
40f687b3
01c12683
00271713
04070713
00270733
00a6d6b3
fcd72823
00400713
00000613
00f74663
40f70733
00271613
00279793
00f80533
00000593
919ed0ef
01012703
008037b3
00f767b3
00f12823
01012783
01412703
000b0413
00f487b3
00ea8733
02f12823
0097b7b3
00f706b3
02d12a23
00f6b6b3
01812783
01573733
00d76733
00fb87b3
00e786b3
02d12c23
00e6b6b3
01c12703
0177b7b3
00d7e7b3
00ec0733
00e787b3
b69ff06f
ffc62583
00062e03
00130313
00a5d5b3
011e1e33
01c5e5b3
00b6a023
00468693
f29ff06f
00008837
00140693
ffe80893
0116f8b3
01412503
01812583
01c12703
03010793
03c10613
14089863
00b566b3
00e6e6b3
0126e6b3
0a041863
00069c63
02912823
03512a23
03712c23
03812e23
bf1ff06f
017ae7b3
0187e7b3
0097e7b3
00079c63
03212823
02a12a23
02b12c23
02e12e23
bcdff06f
009904b3
01550ab3
02912823
0124b4b3
009a87b3
02f12a23
00aabab3
0097b7b3
00faeab3
01758bb3
015b87b3
02f12c23
00bbbbb3
0157b7b3
00fbebb3
01870733
00eb8bb3
000807b7
00fbf7b3
00079663
03712e23
b75ff06f
fff807b7
fff78793
00fbfbb3
03712e23
00100413
b5dff06f
00069e63
02912823
03512a23
03712c23
03812e23
fff80413
b41ff06f
017aeab3
018aeab3
009aeab3
000a9c63
03212823
02a12a23
02b12c23
02e12e23
fd9ff06f
03012e23
02012c23
02012a23
02012823
00060713
00072683
ffc72603
ffc70713
00369693
01d65613
00c6e6b3
00d72223
fee792e3
03012783
00008437
00000993
00379793
02f12823
fff40413
acdff06f
009904b3
01550ab3
02912823
0124b4b3
009a8833
03012a23
00aabab3
00983833
010aeab3
01758bb3
015b8533
02a12c23
00bbbbb3
01553533
00abebb3
01870733
00eb8bb3
03712e23
0007a703
0047a583
00478793
00175713
01f59593
00b76733
fee7ae23
fef612e3
00008737
fff70713
03c12783
00e68a63
0017d793
02f12e23
00068413
a45ff06f
02012e23
02012c23
02012a23
02012823
fe9ff06f
26b05863
01412c03
01812b83
01c12a83
0a0b1263
02412603
02812803
02c12783
010666b3
00f6e6b3
0096e6b3
f0068063
fff58893
04089c63
40990733
40cc06b3
00e935b3
00dc3533
40b686b3
00000593
00e97663
41860633
00163593
00a5e5b3
410b8633
00cbb533
40b60633
00058663
41780833
00183893
40fa87b3
00a8e5b3
40b787b3
00100413
1980006f
000087b7
fff78793
e8f58c63
07400793
0517d063
02012623
02012423
02012223
00100793
10c0006f
000087b7
fff78793
f0f40863
02c12783
000806b7
00d7e7b3
02f12623
07400793
fcb7c6e3
00058893
4058d793
00070613
00000493
00000693
04f69063
01f8f893
00279613
04089463
00300593
00000693
40f585b3
00c70833
00082803
00168693
00470713
ff072e23
fed5d6e3
00400713
40f707b3
06c0006f
00062583
00168693
00460613
00b4e4b3
fb1ff06f
04060693
002686b3
fe06a683
02000813
41180833
010696b3
00d4e4b3
00300693
00c50633
00000313
40f686b3
00460613
0cd34e63
00400713
00269693
40f707b3
04068713
002706b3
02c12703
01175733
fee6a023
00400613
40f60633
00279793
00f50533
00261613
00000593
cc8ed0ef
02012703
009037b3
00f767b3
02f12023
02012703
02412603
40e90733
40cc06b3
00e937b3
00dc35b3
40f686b3
00000793
00e97663
41860633
00163793
02812503
00b7e7b3
00000593
40ab8633
00cbb833
40f60633
00078663
41750533
00153593
02c12783
0105e5b3
40fa87b3
40b787b3
02e12823
00080737
02d12a23
02f12e23
02c12c23
00e7f6b3
fe068a63
fff70713
00e7f7b3
02f12e23
5ac0006f
ffc62583
00062e03
00130313
0115d5b3
010e1e33
01c5e5b3
00b72023
00470713
f01ff06f
02412a83
02812c03
02c12c83
2c058063
408b0733
0a041a63
01412603
01812583
01c12783
00b66533
00f56533
01256533
02051063
02912823
03512a23
03812c23
03912e23
00070413
000b8993
f70ff06f
fff70893
04089c63
41248733
40ca86b3
00e4b533
00dab833
40a686b3
00000513
00e4f663
41560633
00163513
01056533
40bc0633
00cc3833
40a60633
00050663
418585b3
0015b893
40fc87b3
0108e5b3
40b787b3
000b8993
d6dff06f
000087b7
fff78793
f8f700e3
07400793
1f17ce63
00088713
0400006f
000087b7
fff78793
00fb1e63
02912823
03512a23
03812c23
03912e23
000b0413
f61ff06f
01c12783
00080637
00c7e7b3
00f12e23
07400793
1ae7cc63
41f75793
01f7f793
00e787b3
4057d793
00068593
00000413
00000613
04f64663
00078593
0007d463
00000593
01f77893
00279613
04089463
00300593
00000713
40f585b3
00c68533
00052503
00170713
00468693
fea6ae23
fee5d6e3
00400713
40f707b3
08c0006f
0005a503
00160613
00458593
00a46433
fa5ff06f
80000537
01f50513
00a77733
00075863
fff70713
fe076713
00170713
00259593
02000513
40e50533
04058713
002705b3
fd05a703
00c80633
00000313
00a71733
00e46433
00300713
40f70733
00460613
0ce34263
00400693
40f687b3
01c12683
00271713
04070713
00270733
0116d6b3
fcd72823
00400713
00000613
00f74663
40f70733
00271613
00279793
00f80533
00000593
9f0ed0ef
01012703
008037b3
00f767b3
00f12823
01012703
01412603
40e48733
40ca86b3
00e4b7b3
00dab5b3
40f686b3
00000793
00e4f663
41560633
00163793
01812503
00b7e7b3
00000593
40ac0633
00cc3833
40f60633
00078663
41850533
00153593
01c12783
0105e5b3
000b0413
40fc87b3
40b787b3
000b8993
d21ff06f
ffc62583
00062e03
00130313
0115d5b3
00ae1e33
01c5e5b3
00b6a023
00468693
f19ff06f
00012e23
00012c23
00012a23
00100793
f5dff06f
00008537
ffe50713
00140793
00e7f7b3
01812683
01412703
01c12603
1e079063
018ae7b3
00d765b3
0197e7b3
00c5e5b3
0097e7b3
0125e5b3
10041a63
02059463
02912823
03512a23
03812c23
03912e23
000b8993
c8079e63
00000413
00000993
c90ff06f
00079c63
03212823
02e12a23
02d12c23
02c12e23
c78ff06f
409907b3
41570333
00f93533
00673833
40a30533
00000593
00f97463
00133593
0105e5b3
41868833
0106beb3
40b80e33
00000893
00058463
00183893
01d8e8b3
419605b3
411585b3
000808b7
02b12e23
03c12c23
02a12a23
02f12823
0115f8b3
06088063
41248933
40ea8733
0124b7b3
00eabab3
40f70733
00000793
0124f463
00133793
0157eab3
40dc06b3
00dc3c33
00000793
415686b3
000a8463
00183793
40cc8633
0187e7b3
40f60633
02c12e23
02d12c23
02e12a23
03212823
c45ff06f
00a7e7b3
01c7e7b3
00b7e7b3
f0dff06f
03010813
04059e63
02079e63
02a12e23
02012c23
02012a23
02012823
03c10793
0007a703
ffc7a683
ffc78793
00371713
01d6d693
00d76733
00e7a223
fef812e3
881ff06f
02912823
03512a23
03812c23
03912e23
000b8993
fff50413
b48ff06f
00079c63
03212823
02e12a23
02d12c23
02c12e23
fe5ff06f
02a12e23
02012c23
02012a23
02012823
03c10793
0007a703
ffc7a683
ffc78793
00371713
01d6d693
00d76733
00e7a223
fef812e3
815ff06f
409907b3
41570e33
00f93833
01c738b3
410e0833
00000513
00f97463
001e3513
01156533
418688b3
0116bf33
40a88eb3
00000313
00050463
0018b313
01e36333
41960533
40650533
00080337
02a12e23
03d12c23
03012a23
02f12823
00657333
16030663
41248933
40ea8733
0124b7b3
00eabab3
40f70733
00000793
0124f463
001e3793
40dc06b3
0157eab3
00dc3c33
415686b3
000a8463
0018b593
40cc8633
0185e7b3
40f60633
02c12e23
02d12c23
02e12a23
03212823
000b8993
03c12503
12050063
d6dec0ef
ff450493
41f4d793
01f7f793
009787b3
4057d793
01f4f593
40f006b3
12058a63
80000737
01f70713
00e4f733
00075863
fff70713
fe076713
00170713
00269693
02000513
40e50533
03010893
00c68713
00e88733
40d006b3
12e89263
03012703
fff78613
00279793
04078793
002787b3
00b71733
fee7a823
00160613
00261613
00000593
03010513
dedec0ef
2084c263
408487b3
00178793
41f7d513
01f57513
00f50533
03010613
40555513
00060693
00000413
00000713
0ea74463
00050693
00055463
00000693
01f7f813
00251713
0e081263
00300693
00000793
40a686b3
00e605b3
0005a583
00178793
00460613
feb62e23
fef6d6e3
00400793
40a78533
12c0006f
0107e7b3
01d7e7b3
00a7e7b3
c80782e3
ee1ff06f
03812503
00050863
c49ec0ef
02050513
ed9ff06f
03412503
00050863
c35ec0ef
04050513
ec5ff06f
03012503
c25ec0ef
06050513
eb5ff06f
03c10713
00269693
00300613
00d705b3
0005a583
fff60613
ffc70713
00b72223
fef656e3
fff78613
f01ff06f
00072603
ffc72803
00d70333
00b61633
00a85833
01066633
00c32023
ffc70713
ebdff06f
0006a583
00170713
00468693
00b46433
f09ff06f
800005b7
01f58593
00b7f7b3
0007d863
fff78793
fe07e793
00178793
00269693
02000593
40f585b3
04068793
002786b3
ff06a783
00000893
00b797b3
00f46433
03010793
00e78733
00300793
40a787b3
00470713
06f8c263
00400713
40a70533
03c12703
00279793
04078793
002787b3
01075733
fee7a823
00400793
00000613
00a7c663
40a787b3
00279613
03010793
00251513
00a78533
00000593
c25ec0ef
03012703
008037b3
00000413
00f767b3
02f12823
fc5fe06f
ffc72683
00072303
00188893
0106d6b3
00b31333
0066e6b3
00d62023
00460613
f79ff06f
03c12783
fff80737
fff70713
00e7f7b3
40940433
02f12e23
f85fe06f
02012e23
02012c23
02012a23
02012823
ff5fe06f
00052683
00852783
00c52703
00452603
fe010113
00d12023
00f12423
00d12823
00f12c23
00171693
000047b7
00c12223
00e12623
0116d693
ffe78613
00000513
00d65e63
01d78613
01f75893
00d65c63
80000537
fff54513
00a88533
02010113
00008067
01071713
01075713
00010637
06f78793
40d787b3
00c76733
4057d693
00e12e23
01f7f793
04078863
ffe68813
02000513
00269693
40f50533
02068693
00a71533
00000313
00000613
00183813
002686b3
05064463
00030463
00b12823
00261613
02060693
00268633
00f75733
fee62823
0180006f
00269693
02068793
002786b3
ff06a783
00f12823
01012503
f60886e3
40a00533
f65ff06f
ff06a583
00100313
00100613
00f5d5b3
00a5e5b3
fa5ff06f
fc010113
02912a23
02112e23
02812c23
03212823
03312623
00050493
12058063
41f5d793
00b7c433
40f40433
00040513
01f5d913
961ec0ef
05150793
000049b7
01e98993
4057d713
00812823
00012a23
00012c23
00012e23
01f7f793
40a989b3
02078c63
00200693
0cd71663
02000693
40f686b3
00d456b3
00d12e23
fff70613
00271713
02070713
00270733
00f41433
fe872823
0340006f
00300793
40e787b3
00279793
02078793
002787b3
ff07a783
00200613
00f12e23
00200793
00f71663
00812c23
00100613
00160613
00000593
00261613
01010513
9c9ec0ef
00090593
01c12783
00f59413
01346433
00f11623
01012783
00811723
03c12083
00f4a023
01412783
03812403
03012903
00f4a223
01812783
02c12983
00048513
00f4a423
00c12783
00f4a623
03412483
04010113
00008067
00300713
f45ff06f
00012e23
00012c23
00012a23
00012823
00000993
f91ff06f
01465793
00c61713
7ff7f793
fc010113
00c75713
00178693
02812c23
02912a23
03212823
02112e23
03312623
00b12823
00e12a23
00012e23
00012c23
7fe6f693
00050913
00058413
01f65493
08068463
000046b7
c0068693
00d787b3
00475693
00d12e23
01c71713
0045d693
00d76733
01c59413
00e12c23
00812a23
00012823
00f49493
00f4e4b3
01012783
01c12703
00911723
00f92023
01412783
00e11623
03c12083
00f92223
01812783
03812403
03412483
00f92423
00c12783
02c12983
00090513
00f92623
03012903
04010113
00008067
00b76533
0e079263
fa0502e3
06070063
00070513
f58ec0ef
00050993
03198713
40575793
01f77713
40f006b3
04070663
00269693
00c68613
02000513
01010893
40e50533
00c88633
40d006b3
06c89c63
fff78613
00279793
02078793
002787b3
00e41733
fee7a823
0380006f
f00ec0ef
02050993
fa9ff06f
01c10713
00269693
00300613
00d705b3
0005a583
fff60613
ffc70713
00b72223
fef656e3
fff78613
00160613
00261613
00000593
01010513
fc8ec0ef
000047b7
c0c78793
413787b3
eedff06f
00062583
ffc62803
00d60333
00e595b3
00a85833
0105e5b3
00b32023
ffc60613
f69ff06f
000087b7
02050863
01c71793
0045d693
00d7e7b3
00f12c23
00475713
000087b7
01c59413
00f76733
00812a23
00012823
00e12e23
fff78793
e8dff06f
fd010113
00852783
02912223
00c52483
00052683
00452703
00f12423
00f12c23
01049793
0107d793
00d12023
00d12823
00149693
00912623
00f12e23
02112623
02812423
00e12223
00e12a23
0116d693
01f4d493
01010513
01c10793
0007a703
ffc7a603
ffc78793
00371713
01d65613
00c76733
00e7a223
fef512e3
01012583
00008637
00168713
00359593
ffe60613
00b12823
00c77733
1a070663
ffffc737
40070713
00e686b3
7fe00713
1ed74863
06d05463
01812603
01c12783
01412703
01c65513
00479793
00a7e7b3
00f12a23
00471793
00b7e7b3
01c75713
00461613
00f037b3
00c76733
00e7e7b3
01412703
0077f613
1a060a63
00f7f613
00400593
1ab60463
00478613
00f637b3
00f70733
00060793
1940006f
fcc00713
00e6da63
00012a23
00100793
00000693
fc1ff06f
01c12703
00080837
00050593
00e86833
03d00713
40d706b3
01012e23
4056d713
00000613
00000413
0005a883
00160613
00458593
01146433
fec718e3
01f6f693
00271593
02069863
00300613
40e60633
00b78833
00082803
00168693
00478793
ff07ae23
fed656e3
00400793
40e78733
0540006f
02058613
00260633
ff062603
02000313
40d30333
00661633
00c46433
00300613
00b505b3
00000e13
40e60633
00458593
04ce4663
00400793
00261613
40e78733
02060793
00278633
00d85833
ff062823
00400613
40e60633
00271713
00e50533
00261613
00000593
d48ec0ef
01012703
008037b3
00e7e7b3
f0dff06f
ffc5a883
0005ae83
001e0e13
00d8d8b3
006e9eb3
01d8e8b3
0117a023
00478793
f91ff06f
01412603
01812703
01c12503
00c767b3
00a7e7b3
00b7e7b3
00069863
00f037b3
00000713
e89ff06f
0c078663
00471793
01c65613
01c75713
00451513
004006b7
00f66633
00a76733
00d76733
ff867793
7ff00693
e59ff06f
00000713
00000793
7ff00693
00800637
00c77633
00060e63
00168693
7ff00613
08c68263
ff800637
fff60613
00c77733
01d71613
0037d793
00f667b3
7ff00613
00375713
00c69e63
00e7e7b3
00000713
00078863
00080737
00000793
00000493
01469693
7ff00637
00c71713
02c12083
02812403
00c75713
00c6f6b3
01f49493
00e6e6b3
0096e733
00078513
02412483
00070593
03010113
00008067
00000713
f69ff06f
00000713
00000793
f85ff06f
040077b7
6707a503
fffc02b7
81010113
b2028293
7f212023
7d312e23
7d412c23
7d512a23
7d612823
7d912223
7e112623
7e812423
7e912223
7d712623
7d812423
7da12023
7bb12e23
00510133
f54ec0ef
000217b7
a347a803
a307a783
00041737
fffc8b37
00f12c23
000217b7
c00b0b13
a387aa03
a3c7aa83
c7070793
016787b3
02010693
fffbf9b7
39898993
00d78b33
c7070793
04000937
013787b3
01012e23
00090913
20000cb7
00d789b3
00492583
000207b7
6fc78513
c6cec0ef
00400793
00092583
40fca023
00100793
000b0613
40fca023
00098513
00890913
d8ce90ef
16051663
00800793
40fca023
404ca503
408ca583
40cca883
01112a23
950eb0ef
410ca803
01812603
01c12683
00050493
00058413
01012823
a88ea0ef
000207b7
414ca703
00050613
72878513
418ca783
00058693
41ccad83
00e12623
420cad03
00f12423
424cac03
428cab83
bd8ec0ef
01412883
01012803
00088513
00080593
8eceb0ef
00048613
00040693
a34ea0ef
000207b7
00050613
00058693
73c78513
ba4ec0ef
00c12703
00812783
00070513
00078593
8b8eb0ef
000a0613
000a8693
9e1ea0ef
00048613
00040693
9f4ea0ef
000207b7
00050613
00058693
75078513
b64ec0ef
000d8513
000d0593
880eb0ef
000a0613
000a8693
9a9ea0ef
00048613
00040693
9bcea0ef
000207b7
00050613
00058693
76478513
b2cec0ef
000c0513
000b8593
848eb0ef
000a0613
000a8693
971ea0ef
00048613
00040693
984ea0ef
000207b7
00050613
00058693
77878513
af4ec0ef
00a00513
b44ec0ef
040007b7
01878793
e6f914e3
0000006f
00020537
71050513
d4cec0ef
ff1ff06f
00000793
00078863
00008537
c8450513
a19f906f
00008067
04005da8
00020804
04003fc4
00020814
04000018
00020824
e0ffd8ff
464a1000
01004649
c0030002
0000bf03
1100feff
6376614c
312e3835
312e3932
ff003030
004300db
07060608
08080706
08080808
0a090909
09090a0a
0a0a0909
0a0a0a0a
0a0c0c0c
0a0a0a0a
0c0c0a0a
0e0d0c0c
0c0d0d0d
0f0e0e0d
12120f0f
15151111
1f191915
ab00c4ff
03020000
01010101
00000000
00000000
07050600
01020403
00010800
01010103
00000001
00000000
03000000
05010402
00100600
02030102
06020603
04050408
01000103
04000302
31211211
61130541
06227151
b1a13281
23144291
72073362
f052d1c1
43f182e1
b2349253
a224c215
16839363
01001125
02050203
02010604
00010107
02010000
03211100
04124131
22716151
d1819113
32b1a1f0
332342c1
62f1e105
c2524314
00c0ff72
f0000811
01034001
11020022
00110300
0c00daff
02000103
00110311
b201003f
fb284c5c
50acfea5
60feaa4d
f2977ea3
fbf92a0f
417f48c6
cebd806e
b8d72fb4
488bc637
fafa85da
1f0d4d7a
2c706c90
f359e710
553308ad
9dcf1a95
5845896a
433a47a3
225a47f8
568c5c53
2543b188
6a7c0790
dcfad268
5a6cef74
702d7dc2
c698cc0d
06bac958
da00013e
ed622d85
c5318ea4
b37950dd
fabe4601
a2a58c75
aa714410
6cb26f1c
1471f633
47529905
03f2c356
46e671b9
39e4c56a
7c7f79f8
778eaa76
554456e5
338f6578
077cdee3
af28d087
e093b81e
0f00ff06
baa30f2f
60e313af
9ef6b3a5
6d1e9ef1
499d15f0
3fb68173
7ac787bf
08c44ab5
8ce39e1b
593f9e79
a15e8f35
412e0321
d2198823
3ef3783f
db5d017f
e6d44d5b
7ec11ed3
f92a3f67
7cfaea0f
594b8bab
e801982f
6ce44e85
3f17e2cf
ad88de59
45142ddd
2b1f0300
c31c85ed
3100fff2
3524d3f8
b0efe151
35bdf6e9
cb2c5732
c4820d86
3be491fe
5b330586
64159197
a5817405
e080dd00
f1fe8adc
bfdb95da
d407416c
ea5b6937
3fcc4f8d
ca14be49
fd5d2222
c5cde239
7c9e7bbf
9a8cda09
d2ab2f30
431280a4
c7080fa9
ec00ffcb
ec78583c
608ae300
d88243a0
db40fa03
8db36dcb
2d8d1bfc
f2a7508e
ab61a3f3
3b073e98
bd46ee0e
42a74c37
1803c97a
fd5195ce
c3038867
515b5ee6
9c206201
a172911b
1f031675
f1afc0d5
4e793f1e
cc5264f5
1b284070
63bbcf60
4fd4afc0
f94194c2
b16c9764
81b60f19
035ee99f
b1ad71cc
7c6860dd
3cc8377c
69df8ed7
d9af4414
6df7488d
80957862
fac6a6ce
8f7e24b7
9d5579f8
07083eab
6b6e6523
3ee22ffa
e61fc3aa
4e3ab983
0fbc3fde
9a759ef7
45e2a07e
2883d48e
00ffe5dd
8e9c0168
cee5eef6
6331aa89
569f26d1
41e548fc
e5671ec0
8ebac63d
ca328c72
debfe077
a82d4c29
9e989129
cf39c865
858ff470
6c1b3768
2387db41
c2e9fcdf
bfb0149a
44b77fda
2dd74792
0d09437d
b4b11cd8
e800ff72
d909856f
be54a427
2495e12e
e315e182
71746990
884f59a9
d70d34f0
261d1cba
22d75ee1
56e86cd6
386c8c3a
be9178a6
a2e23b57
b11000ff
7f387943
b3e7c121
fe7f61bb
00ff4ca5
a0e1c813
25347695
f94346d7
f2c6a351
ce6a1c91
1955b0ed
dd0ac827
5b3dfb6b
6add0489
9b2fc66e
6e9070f0
dca61f24
c7135f22
a1dba4be
5020504b
6e757262
a909a52e
7d66c0a9
dfed479c
764ff567
c21afe5e
cb1cc012
0243643b
8f5400ff
3d0a3ec3
696fa746
7ba63f7b
976e1b58
12f5df1a
29f5dc34
cfe11854
0c9c4115
bc3f4572
e94ff769
5ab215a9
339dc2d9
50fbafa7
789496ae
4fec7cb3
88693c36
10441b92
83c622db
c4e58f92
e7234dd7
322af9e0
f0e3db4f
6d69c376
63a7da6e
91de3773
0138d4cf
6eae36dc
dd3aac6d
b09cc5bd
a5688ea9
3282b489
189e0a1d
bc23c7ce
cf3c4c56
eaee9e93
c02daed8
933b6d23
fbc98de1
a3f48028
7f993a42
838dfa8a
5b5ddfd8
79dee63e
c6c42762
c5f173e5
3a4e7366
75ddc2e5
e185eb0b
a3c4d53d
1f66e5c9
73a7a441
e8254944
2298d67c
f0ccd5c0
598f21ae
ba4de5c9
fe964d5f
425034ee
a5e9cb6d
e901b0b8
a382d48b
daf73603
7fb60fbd
2b3d48c4
c8a399bf
0058ed20
b3ab8230
63685bb3
018c3182
62146b9a
b7b90235
f499956e
16680b7d
b40203d2
fd46b11e
8182722d
f3753eed
f297cea3
774d952f
2d304a17
0a4d5f91
4d7a84fb
85da3915
9af2c1bd
9c1ee254
3b3f040b
f888d679
8df50755
d5a657e7
ec129852
a02aa215
1c52f155
ec51861b
d77941db
2a3f232c
7cb6dacb
2f275321
eedea7dd
2371cb88
9e449de0
bf7ff7f3
f6bb34f0
465bb77d
dc5a42c6
ed3fdbb1
799af511
666511d6
980d4f27
32307ce4
fd612708
6b2ae458
a31e1686
8d833df3
ee9089a6
e21abf3f
f1381e35
4fe6f139
53f83bf1
a06ea5be
27051b31
cc73c761
dde7e3f1
b989a4b0
ffc08621
efef7800
858ccae5
05a17a48
017889eb
1f890385
ad77d2df
73c29696
3c35629c
e4f3b9f8
56d5f93b
24aeddd6
0bdba37d
977f5fc3
1ed3dc79
271923d1
9f38e009
f4e551d1
f57abc56
0a53a6aa
01786217
fc1c23fa
8facce31
82556c32
c60e7a1c
8c4ffd43
c6c3218f
56aa41b1
1f659756
fad17d22
f5dde24d
c0064abc
1f356ee0
ebbf032e
2db518a6
a701738c
d3fdcb41
52f3908f
c2dd1338
f256e7b7
9ee546b0
9727f019
3452f891
0d3240c4
5c72e2b6
dc5d0e77
2f8badc1
969cea6b
ae3e6c4c
7e87f4d3
e76350d4
fc44c6ee
4d7a0f7e
fc949e24
49109898
9eb1dee1
f08c786a
5a442b3c
21a87451
abefe406
e6e32d3e
7d46ac37
4ec1ea4b
15195e1e
d815ddea
a8318665
fef3950c
b5d6f4a1
48edb021
ed78cd51
3f8f78c8
e2abf3b0
494ef078
368aec24
3e197304
492bf09c
3d2c7dbb
5eb81360
0db8c328
a957acfe
a0b78333
16449d6d
1ee386cf
5330cd59
dde98652
59de99d9
31948f31
c6f00c00
d58eaf06
a1018c6a
e9018c88
ce3b4e5f
b4d2f738
c5b1ecb9
3cf179b2
0af97bb0
fd04deb4
fe9fca59
2a87df3f
29b47a22
475c9b2d
dcf2f400
3e70f764
5fd5c41d
6116328b
d2c0c3c3
fe0abaa5
1c20e9a3
23e8c7e7
2785bbc6
a6c78b9d
5819b838
873c00e1
a0ee2036
aa4f9178
fed1353b
ca977caf
f26cb134
c30789db
5bd355cc
ce5edb0b
24e398e0
38df4e34
e617fa23
8ab18d6c
10cdc6f2
2c3382ea
54793b9c
dcfe6f1c
de51856d
66eaaede
ed1145b0
4fd26e25
d5cfe71c
2b30e0c7
44d25ac5
e60c2208
0441c81a
97a32248
56848545
459445c1
c8d3fc18
f2bb393f
63f7d971
45b0de7a
25268303
54bcfa90
936f1c1f
4daad9de
0601a7dc
95fee191
3cb90362
4042c86b
7d3a0c00
46294583
9ffa3849
33d36477
fb0a3f9e
e03fc965
49887805
dc8f34fe
02a1415d
90e42dd2
3cc9b165
a01fef0f
49a49353
21ea946a
bdb5b321
2d6de449
8f8d5c95
3fabfc13
5dc47abb
4edddb2f
590ab6e8
8f8d10ca
68f62269
c2d4f101
12eaa283
6e65bfdb
b2fb8fda
04fdd5fd
f889cf3c
63edcf50
4f1fcbaf
f79ae9b0
dd00ffb9
d4fe334a
474a4c67
7f6a531f
73b7a580
b5dd1b5d
e264b9a2
f1c0870b
8e1a8f35
b15cc92a
8fb7bb26
1c859fef
c1104378
6580b5eb
8fa4c657
69a1f46e
d6e36c07
db6f28dc
73f1173d
4d368e24
b14885cf
070a0946
d52d6aa5
76f5e9ca
d6c06d6d
6dddc173
56443d16
b0e12b82
975273af
d36c8f43
d375b4d6
2a68a107
8ed67ac8
3cc8677a
894f37a8
7be191d0
8fa17699
a2410f70
3d86c2a3
a5b6fac1
45ae214e
1bebb780
d54caece
f3c6fa0d
a95509ad
af163b84
6c15aa8e
67b88574
8468b3df
1eec46bd
c4f1c522
8c3c96f1
60788e0d
af6ea2f1
b00d806a
8c1c2409
1b506778
e5df4c8e
f64f6840
eb207273
2ec61989
fc1d9a60
8803eb74
81312527
442aceb9
19e670ea
b600891b
926d0c79
bd0d8747
f5aef229
7acaef25
76d30a35
5e1e8739
70128759
60c071df
81914d8e
a36c1cb7
1c35346e
202db603
1bb083f4
c7f1206a
19a2f080
324f9467
1f1082aa
c9001a9b
733846c6
dc66fed3
a3751952
313f9731
c03dc707
d012a57f
492fcb2c
8ee54a9b
de47d940
73f8057f
48d4153e
fe8ff65c
01e4e555
1af7bffb
4a1b6fcd
5ef0c975
67fef058
72deab89
7fbb2b3d
e4e1dfdb
4e03dd28
e99344af
7792711a
c7e0e7c0
eeba7ec1
c875d027
81c94f72
2fa47fb6
d6c49f8f
8967902d
d7e43d27
97124162
3fc3e390
fa3e7f74
b69847d1
0348887f
e342704d
be908371
4e9ef55d
ad12c3b4
827885bc
dea146c5
7b1ee784
e925558a
7b269d3f
c717dd35
33c77d1f
6b52cce1
f382e1db
dd8fa54f
f760b453
ed51cb0d
fa29aba0
737a2db1
f47a4c86
bc808232
a1029232
3d8edafb
8607ee3b
db5bb6f5
b61333eb
12b08097
4524a6b2
b660783f
d48c6d79
d946fd66
79a1112e
d960635d
bbc3ee7c
f7b83695
b2c5e515
4ebc0d64
80381014
73036677
56b58193
1850b99d
e8291075
5f813be6
7d1607a1
59acd56f
359db297
5562b093
bed7bbdb
e66afcfd
a4c731ea
9b15a94b
cf94a11e
f74282ef
4f111567
c9547677
70d5e574
a3500674
81230157
0554f0b1
dd6ca9bc
5946f04e
90419125
6c4232ae
9e14d201
9b22db59
547212fe
00ffbdfe
c8fcafc9
9c3d3fc5
b75c3fd5
5a4c4db7
f25bd255
48555ed7
da0e700c
dabe1a78
37d62ef5
d76e26b5
3a996cf5
c74700ff
d4f8193e
91beed3d
74c1bdd5
112c2f44
2eaec5c6
150802c8
91a83386
8feec792
6c5fa6b2
f6e954f4
cb9b052b
9bdf60f8
593b2e79
88ddfc98
9f8cb3db
1b34890f
48a84dc9
789caf32
aeea6a6f
fb13a654
e3acad6d
262e5146
0f443b9b
dae7a0e5
867be2b0
8e3e8ddc
9c8646cf
511a2386
7c07a30f
3e0f1b28
78ebeb7c
c5e26dad
6a20e3ba
9f4f7227
f5b4ef1a
e11f7e02
d5381348
124ed6aa
929076fb
90d7f213
a0d8ab5d
673e49e6
27ab739d
57aec28f
229a3ec6
a2976340
8ad3ea28
b7502fc9
2cc988b5
16af1aa9
50f80062
a4fd573f
a78f6a2a
8e04af41
ef816dda
00ffc658
4ce511f3
a9d8a2a5
bbb68987
5e9f8186
edd3435e
db0869da
8f05e782
9ef93c20
7ff51455
539a2072
8434cda8
7e78d097
a0baaf86
78e4b66d
b1ce5b52
93d3bad5
4e4ab22c
076057da
ea2e0786
af3dd2db
cf2bc32d
b66b5ee9
a9f19f4f
2837dfae
6ad70191
2609b4c0
b6bf6d4e
bc3aae2d
108d6bc2
6096c359
77152a3d
ccf13cc9
f13d899a
83fe3fd7
215e5faf
65a73dcc
e12de06f
308f47f4
bf687c35
b6fdfedd
d0719f4e
ae6038fa
b18b2b7b
fc1aad80
c88d43d1
78cc3062
2d6a1c8e
f676aa76
9aaba7f4
98aef5fa
981ac107
20ad4c01
d74864ed
c5fa6ebb
f25c9c6e
f466dfa2
9d3971e3
ba7ea5c7
04e8c525
6d6bf7f1
fa94d43a
1e7d66f6
22da58c4
f4869d0f
34fb08f6
4535ed03
27db5aac
aeb8ad80
93248962
0060e89b
575ef3e1
b1065744
fc5982f9
333d47eb
022a5f75
7c9138b5
1fa4f3e8
155da040
5bf82474
9fa13632
6fcb0f70
6a23292a
fc00f718
214ea5b6
f5b8c0e0
de5800ff
153ea275
de5abf9d
ac8eaf66
2e850156
bd23bada
a8e82a52
fa6db865
3e9de455
33eadaf2
90548287
3cee947f
fba6da88
89319780
4dd02a23
38657418
04b98c52
1c54011e
0038c113
ea78a05a
759ffd4d
e6edae89
da7a12e9
e7da3224
1fd5e792
4675927e
a87b320f
34a85317
8c8508ba
b3cfedb1
846cd459
8ea3f24e
230192cc
f1f7910b
b0f439fd
9d73f06d
174552e8
4a231753
78ae4a67
573f050f
f741aa1d
b2b7b10d
acbf4694
9ca88d60
bf750e46
2a9e3f8e
2299b83f
063a28ca
95e339c8
96a1ac35
4d7e0975
63448f2e
3cca7f7c
a8577d4f
e3ea132f
75aeeff1
c9b15b24
f08fbf63
0d6ca4aa
3f780067
381e3ea7
a9d901a3
d3d1ee2e
39d49532
ce3c4a0d
7acb031b
6dd47fc5
154b0ccc
8d626474
090e38e9
66f8f1d8
a53ef5b0
495cfad8
58cdfda8
8d7fb55f
cbd14c0e
b9299df2
1e4fa2c6
a377fa5b
0aaab1da
ea1f7584
89fe7ac1
8b430f02
ecbad4d5
13c24597
86233914
b2ed8eed
90c27e4f
e7237bcf
ee5ce842
7b72eac4
c23ddbc9
9d95b9aa
1ca4cfc8
aeaeee05
c6db4a15
b15c289b
e48ea9e5
dd4257f9
7c40a0b4
b21497fb
7f972449
338f654e
caa7f2cb
9f9cfa0e
755adfe1
fa98503f
e314289a
276eea6c
1dbb390a
3471c0f1
abaccaa8
8d14701e
97ab71fc
94dbb5c6
ba1d22ed
a8a80de8
ee18b90c
e91d791c
d4303fb0
5cf6641a
8da4ba3c
7f29a807
6b042b9b
a8bf99f7
6972eef8
a5fdb7cf
b49600ff
def19eb6
2bed420b
25f31b48
287bc52c
a862f190
03d8b9a4
284b745c
b9205926
29752b66
35210079
85285824
6c09e18e
02c0719c
746a4fa5
7109a3c8
91405270
1d401481
a063a810
172ce563
e97b208f
110a3777
1c23a1e0
96ac6e87
5519856d
e8b1c940
f08fde5e
f8c1a3f0
fc189f5e
ed38559b
cef9fd34
e9bb99c5
084085dc
005e8406
1fd81d70
78cb56e9
b2ca31a2
3bc8c176
2a06ee9c
a9318020
504ed467
bf3b1c32
0ce0d911
538eac62
df00ff26
18628d97
de8ea9d7
cecbb31c
2fb22ab5
343e63a4
f470e4e1
3303d509
4ee20010
b72ea1d8
d48640fb
414d07cb
eb603c77
be429c90
84bc713a
e97b7a77
b8a1dded
6288d585
f87083c3
3a8a1a7f
97e9a8c5
2a18ae4e
e06eba93
398e8f7e
7acbe3a1
069256f1
d0c23647
7b329e20
e59d3aae
d43debec
d4fa7ce6
7d23d0e7
a030aab0
d7e2740e
87cf58a4
06c42e65
f0c7b120
b85b0ba1
8905f6f5
38d13259
c9c84123
97d7b903
277adf88
0b4afde9
24ce3508
57018370
fc86638b
d54937ab
5832996e
41902920
e8601463
1a45a058
0355b699
db872799
fdbdf751
a45f8ef4
648f89f4
8857b732
c578db71
ff110e0b
9b0f5300
dffd87ca
b6ee9bef
fb5f9c4d
9863354b
0ef32723
2d6edd7f
e384c2e5
9ab66daf
70e2b506
dc5f311c
34a584f9
77ed1203
eeac0acf
71b8ae40
6d4d60af
f0aaf2a8
28ae670e
4789948b
065d4a9d
e3ec6ccd
064c8d41
db1be87c
e0e226f6
9a1b3636
7d4c3a92
2a3fd9a4
e92675fd
f7dc2758
4a84ed74
73b3c3b9
0284166f
e35d2bad
35ceab6d
445da61b
35ae0657
aee71559
abf58339
1c9d47e7
ad8016fa
be5800ff
fed17b74
c95da145
e7161899
807b0d95
35515b7e
e4837b0d
3dc4186a
4fc7054e
35f3d6fa
50b531a6
ce5bf3e3
b52ac6b4
5f9cc264
0ad15540
7f9b56ac
b16dab4b
f8c8301f
5986628e
468ad003
b7e73132
fb63741e
3a48b83e
f9f141ec
e7124bd1
0f04309b
84669c8e
d99546bb
4eec72e4
feb9134b
59ab56f9
3996b6e4
46326d62
1047e8ea
db0f72ca
945e5543
881c496b
3eb49f67
1dcbd1a4
9d127b9c
ec7da4a4
1beda793
92e45191
7e323ceb
765fa2e8
b53a48f5
edb017cc
f6d1d624
d749f3d1
b17dc32a
43e5189e
512fa26c
7fe23120
ad789787
916af5b7
9066daa6
65d2dd2b
56ae714b
ed0ce404
f7f72485
d5b17ed2
cd7eb057
e91198d5
7c1e1ccf
d5b99e6a
95a64c20
813c8590
0f204ffb
dcdc097d
437b70cc
503a83f9
0f39219d
f66d57e7
23a370c5
c66d6ebe
8a945be8
9b9e2cd3
c934a1ee
baefcea9
791c887e
a6e8d2f8
7072df68
7e00ff78
da8dd475
4ac74d2c
de07d284
15f3f104
ce51e753
d5f93832
804840e8
2a6a3d1f
39f72e33
b75ac30b
a0452bda
afd68c49
7164b4cf
0e4fa6c8
86468d75
46c6594d
7670864f
97de1af8
6b714770
55b09134
a71f7370
91d7ab2b
6dc49383
78349dca
2a3ad66a
cf874be3
cff31871
6c0fa3f0
e3594afb
1be1f28e
76f4bf5c
fe5f7adf
3c751fd7
bbcac733
49d43ee8
b9ba256f
cdb1764d
ea1cdaa6
d71d4bfc
d536c6bc
77a976e2
0dac58a4
e1266dae
84ed18f0
78d4fe41
d9977ed8
24b7ee51
0f072d1f
8ffc5fc9
b66da3db
ffb198a7
b33fe500
bd2d69fa
684e17bb
660994a4
c3ca3166
40596305
df18621a
b29f3146
1c962d8e
30a43112
5f3e875d
9cba58e3
a25d0c2b
9d2a71ae
cee377b9
6be9bcb4
c9604368
7878fb26
facffa9e
57230ed0
524356a7
350fe774
83248dd4
b69fd303
8c6596bd
49b59508
b8771fcf
2e09d6f7
1c4a4f9e
57e59f78
1ea343db
f195a179
549bcaea
5b7c7a95
1575283b
1823ea2d
698af7cf
1e9e82d9
04d79655
504cb10d
13d1770c
e9e24583
ef946536
8b3a8fbf
d160fb3d
6a3cb0be
ff304c64
f7024a00
66bb96fd
fd27cb61
c1a72f6b
b0bd2a23
300751a9
a66babe0
b1311e49
c1a3d647
f1b8e3f9
bfd90ba3
5b1600ff
63a0ce88
80dabd0c
4ea0b7fa
c25b9ba5
00ff6cc3
3ddd4503
eeb7cfc5
e78cfee2
9053fe6c
470cecc3
00d59cc2
00ff40e4
14923436
062cf1a4
1223cd60
85af1f0f
f96aa374
f03987d0
157d39fa
47e3c8d0
2e6130c8
4cab3cb7
c0ab8009
3bcaacb9
ef343e49
367ed9a3
54c635f6
16ab3c10
52e58a74
035101fc
fbed6996
2b5ac30f
2826d763
c32fd2b6
e64e3c46
82dbd8b1
637a80e8
d4189d02
afc55ced
dee58952
7000e994
76805bfe
c15a573b
09936ae0
65155ce5
a7d7a3ac
ac09ae39
7d2fabdd
7880f875
fcd25eed
fde08f0b
e7d1f962
e117f945
edb81040
e83f7a17
50f9a29b
46e8642f
bfa1bc05
a8ad7e70
fe3a8796
a1913f34
dc8c5e8c
5feb2773
bd47b4ce
aff59767
3ca6d5fb
ac548d63
b08b9398
1955f155
a7bf351e
287d4dda
1b69048a
9d209d04
63b3382a
85341e80
c6c80ebe
e284e97b
c5d8a5d7
5e69297d
22882a43
8274255d
b3da5c17
4edd311b
ebadb093
9c4b8fd1
e55172c7
37c85245
04675808
1c5000ff
a88e2a7c
4e5a38bd
0ee56ab7
ba9c1d96
7ee74a19
b8ef4a05
55418a61
07d4c40c
06093eaa
ddb47a3e
d5c7a81f
dad1f0d7
83e16cc5
f0492afe
578620a3
9ba79163
37306e33
fa567dac
1995162b
11884696
8e9521e8
056e69e0
4a118f39
4da7faaf
2c0e37e9
e0527920
78ced006
18554010
3e69bfd4
e29aa114
a26fcfe5
5c160015
a7937182
283ff151
9d75351e
206594aa
4f9c07a5
6eeeb8dc
ea041342
1d309c50
fc150f72
f059c88c
02869d64
f7ab008c
908ce340
8b6ace3b
148830b5
920126e3
b74d8d39
4cad37da
05b7b484
0a764477
6563424e
c29a7efa
3c8665ee
e7acc9ee
39d95299
1af93bf2
211200e9
2449d4f3
4449f9e6
a2bed263
e0c7733e
aaf17939
ef07e786
22d62a7c
9091831b
57778cad
ce18db53
be89eab1
3cc65d57
aff3810f
d9d5c73c
96db93d9
a44b6d18
1feaf11d
fa4d9152
6a1d4947
8b7643eb
2b336869
f50754f2
24ef8c71
34fe9dad
4e5cdcae
6720dbd1
c0623a77
1a98ccc9
3c1e714f
97f6642a
b7b0e3b7
285e3a55
95877698
27dee7d5
c387e36d
759f0a87
244ccb7f
19f488f8
c5a2839f
0f954a9d
1b9efa08
25f46f2f
17635685
20002367
84b78087
00ffb68d
f11bc388
759a781c
58bce8d8
6a9c1e53
69fcfc3d
31f6aaa5
76eaed34
78e90fce
f75e97d0
15b7bf4d
df323dd6
ba8393cb
3f83a7c0
9f2a1e8b
8446b513
f8c84f60
c85c4997
01fe7d19
a59ef590
1de2d36f
c79564a6
b6c605a6
65e70cc7
a86df35c
75aeeb26
2d492333
f2f358b0
f403ab27
f838899b
e7355077
3c3325bd
ac2ccd8c
25c7ce72
87c7f08f
be56550c
3c93eaee
93b485fd
45e58beb
174fa72d
51780220
baaa2e4a
a55a3d61
291e9176
402e4157
8c5df7b3
c66c168e
6d8a4a7f
23eeedae
f98a0c0f
590c35f0
8c7a4875
b2532e9a
b865c072
cc970f0c
2afa1e9f
646c4ce9
3ce96dc4
ce122a47
cf100a83
0695f968
b54dee7e
2fc7c1b8
312e603a
e72edd42
6adf75b5
636ed46d
897bb7b1
5d44639d
69fa38c9
1e45a290
b705405c
45c900ff
22f2d408
01bb3380
7d82cec3
9fdeeedd
1bc13224
f283a4ac
1e35ef9f
f0de83fb
c7d1ccdd
a507ceda
ce4d3840
1a1ac7d9
c753dc97
b16e0323
5c96fe36
14e61f30
9816375d
18cd43d3
5448cb4d
8767afea
4df34aac
f10da492
3e7b14b5
b0373c41
ab59f313
fe65810f
7b7b2954
f90990f8
c63fd08f
bd913d89
daf5afc3
e463bf48
002d2251
4c124344
2c9999dd
323dee7a
9dba813a
3c187324
bfb2c647
9fe97ca5
d4fd4f55
9c0d7384
e9faf178
072ca75c
0654741a
7544fe25
dc215b7d
a3bd8ee2
721a1166
0e9ae137
50155cb7
28154932
c63e8bf4
ddc018d6
ba812680
fb39265c
2a916d33
9bee1b9e
9ef5981e
cd6ebd2d
05228056
5475aff0
3e8aec12
72bee2c3
5ef3aa08
9017b466
aa0664f8
1357b378
b215165e
ed36c6f1
52e7c9f9
843e4147
07caa8f2
a9f3d4fc
e537a02f
700f95a7
71b46630
86da5864
87bec0fd
501b75a2
a107b8f7
1603a8bc
edc6cde9
9d37e71f
beda235e
9db7d66f
92544168
da9907d0
c291b738
cc0f90ed
cd73747f
cf9df63c
daf58a50
bcf4ddda
619ca10c
1be8ec0b
00125870
59ef1cf4
dca7c396
9bb8bbb8
194b244b
942b978d
8daa541a
818d2bdb
3dd59ce3
6d0fdd43
99684732
e4271728
53f4a751
98211ee5
994fdbd3
9e318944
5316570c
cb098c3a
fe7be412
2a5d049d
7577b54e
ad619105
bb5959d2
b8453c67
89d90990
7e0749db
750c1507
cbbd74cf
f83604cd
ce129c77
06aa6249
0fe02814
ad97f576
acef82fb
ed46665d
460c1888
e5033416
a30a178d
8d4f3c6e
b52a6d73
ed9969b9
b7235d24
21e62f8c
936c00ff
6d0356ea
5d9bd540
55551382
5f3f4d5c
dddd2557
bc424ac5
e763c53c
d9f5b536
cbb56d9d
fbb74b12
1da4bf7a
551e0fcb
a923c55b
ea03905c
3ceb9124
72649ed8
a3ceab1c
831af1a3
0408ecb3
237d861d
dc769224
dbb4ce93
84267183
dac91c60
91f5e32a
7c9525b9
6e157258
99e53098
c2c25e77
724eebda
04400082
fc7c2767
2367a477
79b99d63
d3aea2f1
ab140db4
35fac82a
7d17a046
8c41841e
7b3e48b6
ba1a0a1f
00ff9a1f
a511f520
e3e04232
78fbce48
8850a7f3
38935f6a
741c8694
51debf2e
35c0e9a7
6322c9ca
b6e3304b
5738fb76
f4a2c714
b1d7eab6
dd940ec0
89e87fe5
03fe6677
04a586be
af024e02
00b29252
63cfb2c4
99ab6b74
d058b821
7634334b
4ce9b3e5
1cc1657e
a7904100
e9666a1c
a3485956
24864445
134ba3d2
49727780
9d3ba71e
3ab60fa9
b1cc887e
58754529
a5605c62
f1c170b2
00fff190
3fee691a
adb72770
5706d2d6
8e7399bf
09cf0822
b89f7818
b5138fa7
aa797573
6300502b
0d7d90ed
d316583e
bec48753
18eec9fd
d6666cba
e95c4bd7
20441cc0
e3b800ff
bfba1f9b
3d45b513
5f5ca44b
69eb922c
a3b6640b
4b3c7696
e634391e
793933db
6a33bb18
13cb6d76
224e93c4
3e3dd4b2
52e9a674
668065a4
c104dc4e
6d5ce2ac
65bbb717
9528b1d2
82d99873
1eb70dea
a4da084c
b6efd93f
d748a79b
41236e17
ed208909
3996b354
517e4a32
6fa06ca4
452f59bd
cc096332
ac668e9c
8848a283
1491b517
91c04e0e
a2416e8c
32b0f2a6
8853edd0
dd7d78a1
ff1e6cd1
d016f100
66ba12a2
cecc8fc2
cbb0e9ca
30a5882f
0cb891ac
f9071877
ebe87cd1
c5682f1b
2c9fdd71
6a8fa4f1
0b747e13
77cf38d5
4044b445
68ed4b86
2e32137f
b0c69178
dc75d3fe
d64f2fdc
f1b142d1
874c3a55
438ed538
68dfd6f8
3ef25248
f0bea7e6
485d32b2
aad688e1
e3f61c48
e89fb246
c5d43192
27c1fb7f
d8069702
f1f35efb
8abd4624
39f2d2b8
2323cd4e
649ba70d
aaf0ef70
5204e17d
168c2edd
c6a5c655
e8fc1d49
4959a8c3
fed6311b
23968ead
cd0b856f
66b1b4d3
b13810cb
c6a7fd24
4325cfb7
b6951822
a0024909
2f1bb3b0
3d8c261e
56eae897
3a70fdeb
43b359fc
6f7e11f7
71d2bec1
74b07d4f
586e8b75
28fdab4f
8fa45eeb
e9b43d57
75f3ee58
704fb488
228f8231
3e8ef98f
faf2d08c
6fd1f8e4
beb053bb
2819dbba
c3d4efd8
758ba1e9
cbb7efd2
41a6f3b0
45b9b5f0
f6dbe716
40be887f
ee39c041
185ba5da
a3e4d9f2
a3bd8202
62da886d
f628e037
0f113dce
dca1de16
8ae352af
d2e9f63a
46afd681
9af8ca6b
7f65a7fa
ec2b9c57
bfd624d7
25d5183f
3da6a6ab
7a4ba337
ef842041
092a5ee7
2ef64b12
35bf851a
f64eea7c
e1d3eaef
7ebb5d51
a5c6676a
a9fe6e2f
c8ed153e
3a83b5c1
1f6a4899
daf2c7eb
b91e529e
4d953ff2
71732a9b
6fce1ffb
4403dd3a
f7335830
bb7da403
61c5f093
a5778d40
32b614ce
e1330f78
111cdf9a
30f9fac5
101a8173
3eeaf758
d5fbbd80
8f88497a
17032976
8257d7cd
b455fec8
75d9282d
1c070899
f67b90f3
f55f0ccd
2ba1f92b
58886627
638962e5
4800ff4c
f33bc9c0
b7a6ee39
52d70c57
40916ec1
bff3d4a3
803442aa
32865b70
2705d200
437037ea
994f00ff
37ac7e14
af0c5c0d
4a8f58e2
1b5d338f
71028009
1e08a422
d4ea1bce
4003cc4c
9bbdc2f1
cb032a20
b7f75195
1c72c4fb
9abd6885
c4a99018
b1d420b2
1b5de981
6181db65
6395c3e1
9225495b
bc0a6927
77be038e
776c7607
93dd8122
6dd5d38a
0ed346b5
477d5938
1b6346e7
150ecfed
b66835be
855c8252
91275a52
72ec72e4
dbd6e4c4
1240b06b
3d66bfa2
07279d24
1f8c7190
b0a2fd0c
afd5b691
a99b59a7
1c801254
271859e3
f838bc7d
90a094d0
c90f6954
59812a0a
48aa976d
221024b3
f9ab6c27
d2b8b9ec
4609bacb
ce953130
ebbdbee7
582b36fd
08625896
bcabaf84
fc1d948c
bd5578ce
3211a63f
f4228e7a
c6e51b99
0cb7c072
89de802f
fd36acfa
2eec582e
5f59dcc2
4f2c6544
5930eaca
959fee1f
2ea9f0f6
0c5a096e
e65c4695
a675764c
025381c7
b8e4e373
65efa4c2
22580674
bd67e188
fe1b4922
14eeba1d
cf65dcf3
426750c0
75dfd1e9
a11a1021
3f776746
78f890f0
53e3c3b6
e1adb587
eabab6b7
88617a57
38c7fc29
768be148
0318f039
6eaf18bf
da9415ee
a05fd519
2d8f6cd7
a072b82a
abaf97fd
694fcb75
95baa674
82484843
d79fdcd2
3cd2a74f
7997387b
1635f10f
d4717b41
e6ee9267
31d32c43
9fcc6377
0038000f
c56a0336
b773dfee
53dc7abb
84b36420
3b22ad98
e6cf2562
2bcfce15
b0e14d0d
c2f45ee5
79850257
ea13101a
b556b7cd
26837395
9a116cb4
6c90b224
5b0c850f
2d4f313e
c9541b64
0a445f30
95c24832
677cbcda
17242b86
e170a00a
14d9bc56
2963545d
605df282
a282bbd2
164cdeb6
6adcdc91
925143e7
ef0d08dc
780ba4b6
146a3b87
81c1ee75
20ef8304
0a073c1c
d82c7a8d
7a237799
fce8fa92
b8b64347
7794111c
dacfe5e3
9ba99d6a
73150737
b45d84ee
372e65ae
38098aea
55ee87da
cb937244
f59fa26f
9ea1b913
cc8230ad
55ab8193
d44d5504
62322c61
4fe4cd0c
a9fa76da
1d6d43a7
4fcfd366
a4f30fda
ee6c3f90
c9c3d5df
d234fe76
aacb4ec6
f1e4b85a
50aab29f
bef64fd3
ff994c7a
fd6d7000
c73211f3
8232c830
3f19ce87
22862288
f9b0938c
8db66fc8
7b01eb7d
59c9f822
a2dd1d81
1c9afe8d
e2c636e9
011c14f6
9700ff00
6e71a115
53b79778
67986337
b1cf0a9d
6e3c82b5
a2f113c0
15403a8d
82c5a783
5354d936
3271ae16
10589767
9c6bd621
22b946d7
245ffab5
35be26d7
f2343164
8edd282a
3d3fd82b
35a723bd
3a88a1ec
da68fb01
42dd5608
d353c5a8
05ce966c
dc8a6f00
2bb63391
b8f17e9f
a03618a8
e0947f15
9da7da43
04dd9e4a
eba89944
651e44a7
f42635ee
571ad385
e8587143
076960fd
1f297cab
795bfd5e
a4c9a453
5b7e78dd
a9ac5479
8448d171
c77364cc
7e924164
265c053c
55e8ebc6
ef76dcce
58df13cf
f377dae6
66c270ad
a00ac947
ed82e76e
fface2fd
2d1fcb00
699e971b
60a4e10e
31247135
18f240f9
8d6157ac
fc3482d0
6b1c73c6
7d8ccdb6
2b3c99a7
9fa53ca3
26802493
63d8789e
6692679d
26cde4e9
1090ba97
120afea3
c3a63f77
b1d515ec
e92e1f40
c2ee9e04
6fc75ee0
99486392
90660701
f76c162b
5b31fb96
59dc8067
0020d7f4
84942dcd
81d2d2e3
7af39fa4
cb52f794
8ca48d76
765b7ee4
d5e62383
783e799d
5ac556a7
d57db617
f056b7d3
45bbdd92
b7a0dfd3
3132559d
0b8acd62
41c8d676
78aba4d4
27a70d29
d2df7ac7
b8b7b7e7
c8ca3ad3
32d9d51f
f9a9ba2b
3cc0b054
b583e377
68b2be6a
01ee84fa
29e62f29
0c51075e
e0fb1dc3
b4e0de55
1e489eb3
8cc93ec6
820ddb6b
971a1702
b925f018
b1b8a4e6
0633cbaf
caee326a
429d1094
9b3d9729
b7b2fa38
431b9c4c
ebcaba15
2249c31d
d96f2393
665013ca
95ce00d2
8ba1713b
dfaeb99b
42309056
1a671ac5
09d2c088
3ad34534
8659cf45
2dca0a13
a01e93e3
c481387f
8927639c
a21838c1
d3b13d19
dc313cfa
b6bb2e5c
e480923f
53668c26
0380cb91
1b9caa1e
49a00a76
e5f5f4c4
e4e5a69c
eb324da6
4f74dbe8
63634364
27998d18
5dda5e74
c4ec539b
809dea7e
ebfbdea4
0ed85bb1
d20c2e8e
71248900
0a358e31
43646943
750224b9
9bca9313
f6e7755f
e46944f7
e2edb59c
5f85b015
5507d368
0371a0dc
9bd90682
2b4bd4c8
cb2b75c9
2bc93323
593c6797
994f729b
478db2ad
32c954cc
0f6075fd
8e02312d
00ff9fee
880f6c51
2c899afa
9ff85780
86ac87ae
783f988b
d2be1d51
dca579b7
fdb56f99
18e796b7
1f5b9cde
e101470a
85df6d4d
c129fa42
152346b8
2fc559a3
b5e24c8e
4ce3c8a1
d457f30b
141fd59d
6dedaead
21666284
3603869f
221ac04f
1090249a
9235fd79
3892922e
1b763c03
1787751e
61c7a3ef
0a4c127b
3f7eae1c
5ba4c611
ed8db4be
c928c2ef
9623e873
52f99ce0
5b695f2b
c2057845
604d0199
1e2e4f67
abef1a9c
8d285aaa
18854217
3d0ac051
56daaea4
30442466
942e525d
813a18a7
c85f8cc9
81c6a74f
37d4db7d
b73c645b
a2f15fee
b676a99e
708ca4fd
e093a4a8
1746bd31
33772f97
935cdcca
f0010fe4
bda55d14
f7939c4a
696fef73
be8a914e
e7805dcf
c959bfe0
6260abfa
00ff2b93
53853f46
9f8c9864
074e1fd0
3e4a57d5
c1befd6e
32eb94fe
0891c0b2
eb42ae1e
271db74a
2b5c0738
8f00ff27
96d99314
5692a745
e7032f1b
db9b06fe
858ef8cb
0b71fc6c
3f0ddfc6
b33d5be3
315bf865
f563b991
ab7b2aec
92436dd3
2d354ae9
862ce12a
efa134dd
86af09ab
727507ca
facb0d68
9a79cdbc
f2f1bcfa
acb6ef69
0819b3c4
235278f9
8bdb9e46
3b3eb845
d32a77d0
336cf56c
0067426f
bb780b53
5d759e31
1af559ac
b75853d9
fd968bfc
778ff0d9
e4a527f9
2675be4c
6b4c8074
1e49b751
4caa7cb0
4f68e4e8
b2fbbe2a
0aca0dd6
e587d74f
553e9537
59755da4
1e727ca2
b9e36d20
469380a9
bc199744
2ad32d6d
90c7d5f1
02eec91c
43a334b5
e29860ac
60de6f46
03fe763e
34777995
0c869670
e9fcb9b3
3c117c3c
b9267d14
dac17fbc
32c3193c
5be05366
56219f82
b3235524
1e058c12
953b6aec
6590d94e
9c7342e3
0b39887a
91268ee3
49d4f9b6
cec98d24
f7ad493c
479148b0
3a357026
707207a8
24723b01
189e15fd
d80c457b
fdc164d2
fc5b30d0
9175cdb9
d4a57c80
468e61bb
7d803288
a5461f47
b0ad88fa
6eb432cd
19e11daa
b9bc9f31
94faa3e2
b6c2631c
ba6d6e43
2fa19418
3fbd89f8
199071fd
7a673e87
c32615a9
1f2ef22e
8fc2a563
0ec431bc
c694a278
dbe6da1d
f8044b5b
34dc509d
9b186631
158aa909
85c01311
46e2d338
dbf79a38
aa97dede
2c5e32bc
94a3fdb6
9d6f3c88
0fcf6763
ca23f049
2541dbb2
5a85caf4
2ab32707
633254aa
19e03850
a4e6f8b9
c392825e
81e3d377
4619ca43
512a5f89
b618587f
a87260c0
d0098bb7
41ad5440
dd693e26
56b6b6d9
01422415
d7c29650
5a6d8fa0
8c26af99
12651b43
1b799d2c
4cbd5d04
0a5d1f48
7df10b75
ea54d72d
b69d4507
6a9c1a33
9056f63b
89e76e9e
a8dcd4f0
7257dc97
4eee927b
2c2cf2c3
1e60fecb
69e91480
d3c78e07
51d41c9f
45708fee
9515717f
b34e479e
fcf2d92d
ee61e444
2a3fc75f
e3f08267
d5454240
18a18a94
960d4f9e
680284a2
0f3860b5
9f52d705
5eddddac
a583325d
928d714c
86649338
bb8ae425
d63bf101
c7488648
11673f26
98b82c54
9faec093
2060ab81
e2c37e65
4f4c51b5
33304761
bed44bec
fdf1889b
a9dd7e6a
43eb6fe4
26f083dd
a27ab390
e300ff6e
93a24c91
a3feb9d4
892ed0f5
55f6cc1e
c092dd07
0c610adb
c776a598
6cb45620
8abe881a
d7926a4b
8158f93f
8e0cda29
538d8d3b
deb1e60b
2577dbf4
be7330bb
8af6cd46
3149efce
bf6df748
139c31f2
6b8d8f22
7676ebb6
abcdaeec
f56de01b
70569cd0
1d096eab
e52972ec
12e9459f
16126728
3e60ddc7
682a22ba
24cdbb47
66a9078c
a5cbfb32
d6965bb9
834e838e
1c390422
c337604b
b98ea1e9
e66b3bee
2ee7f08f
470eea4e
e5e5f576
7d4b459f
5de6c031
79831d86
92bd1d9a
4c0b9d0e
9c141ad8
0e78c001
52cb68f2
894a89c8
0acb00ff
88758b92
63a0498e
18eaeefe
f556b454
fbcb7548
273eeca0
8b2a14e8
1f3f80a9
2eabeaaf
e6fa5e2e
d9e2e449
0507e06e
566dc01d
2497c75b
1fc7faf0
4542adaa
89737a9b
2de6cb3d
acc2757e
d96007a6
8e10aedb
57b8fae5
710fec52
5b5de3df
fa0765a9
74c5ea9f
bc975057
a522ec67
2c3c9ecd
77fea0bf
89c40944
46e63f59
ec8aca1f
41e3ece2
bfd0f4e5
b55dd7b2
2abb9fc2
a377fb30
3e2ed428
f2e33e15
9b2eeb48
909edb5f
35b826ec
4871aed9
b3aff9fc
af99575e
e6fefc10
fcf6452a
dc41b719
e44d3a2a
eb43fa41
40a167a9
c41bd112
9584fb54
6b594fe8
b55d7e71
2cd9601f
bd02177a
d65e75c5
f2f97084
f42400ff
394488c8
7d4845e2
1e10ce15
5cfa8fea
4046d59a
e83f8a00
543ee5c3
f525f34b
327b44ed
1e52db60
e56dbcbf
5ed2944e
f2a6fabb
2e4e37a0
3e968939
4ee496a1
db58fd33
529da5e9
604c9969
6cd9ce82
fbe758ee
799b98de
11e42eae
5d50b923
086da9b4
1cdb25a3
d2240e14
c62ca10e
6455b3e3
38cc0e24
e7ab29c1
1d67dcf0
a7dbd0d5
e5408752
47122adc
75f12826
dbd1805b
183b06c4
4b2ef3c8
d4a9b21f
c6d122c8
fe69c328
7c367fad
edf4dbeb
e9839026
c727146c
b3a29f86
d46585bc
ff402137
ae889700
8f864f8a
ced4a99e
69111a2e
051656d3
c76581a3
762951fc
0ccf3692
b193c2ea
e5056be0
6d3c71a4
50159a14
27a348ba
01947a4b
c31138e2
eda21a3b
b7961665
f62a3331
117c8070
9f8f8d94
7267d52a
aa438f64
30352eb3
4e9f391c
e7727cc3
ea54b38d
0f948606
775caf22
e1052c6d
d0c0305c
67cb2137
71185eb4
c1e9e0c4
dacf28c6
aaf302b7
86d02413
d2d0b854
13680fb6
f549ba0a
08d27690
415b0acd
4cf94d0c
1ccd1caf
6b1d2380
08569fa0
074982f4
ff71778d
d7e99100
9f62cd93
aeca0a98
9c415c13
245b196e
c3cb6c1c
5bd4d850
92cc2ba4
1e241d24
aa8b1f23
43b780d2
e139825a
f742fbf5
fe17475a
8d48a60f
d500ff12
da81c55c
c6d8ed3a
73cd6e57
4e4c1dbf
32441bf5
c4dd55de
48f9e4a1
3b69f454
df921337
fb494ea4
d455ab2b
d5b6cae7
c0eceda4
96cc49e2
bbddac05
107c703d
fdeeb735
8dba669b
ef19b0b4
f397f55a
3f15fd26
3be4aaca
a7f5afbe
b30f7bc4
efa51ef6
727bcc66
d8045ae1
3f08bc01
7c225803
3c3c1e8c
30cef4ea
54fe8847
6e312215
beb1250b
e24e3042
6c30479a
763bd060
fc912ca0
a6f188c3
c64d3d56
8e54403b
58aea939
d565a0a6
55fc736b
3960cdea
cbec6cc5
a7fd508c
93638b55
4ee51ff6
7294baed
7d2afa72
4aea6224
53bbc0c1
6a8434a6
00ff6a1c
d5200bfc
011e38da
bbb5318d
370e5047
97446be0
0a7f8708
d2cb8170
16e0095a
518f42aa
7e92cde2
c9bd8f9a
97c44dd4
45f42911
23df33a6
50fe5b36
7db4fd34
b5d5aed5
38652395
af8a2ac7
7282a40f
cf91465e
d1e4f6d5
7c05c9f6
1cfd7cc4
9810b57b
af7e7ee6
c6960b24
c8ece338
388dd1ad
99cf90db
dab3ca3f
bd7f5b2e
2fb5b29f
603fc7fd
9aaeaac0
0188edb8
951fb6b2
f563f109
9f0fe88a
55f571f7
17430c91
57a41f9b
d29f6dc0
900af71f
61405d9c
3dcbf4db
8b173d8e
078c86fb
e2c0c3cc
e9953d84
fcf2403d
4493f6b1
8e23d44d
42e35346
cc0e55bb
de3da2a9
d6ec6bf2
fe8dbb55
072458f5
2fb11481
5bd5f625
54b5f81a
d20f5bcd
68268bec
eb63fdf1
21a6a3a9
fe41384b
3d54f591
3737e2d1
f53746f0
d41bf083
120918d3
551f058f
4eaa510d
a31b2c49
5fe548e0
737cdd67
89036b5c
48bb65aa
b550dcc1
94cee1c8
5f824629
399f4ee4
38ce208c
f9ed9354
bae3aac3
36a049a3
de7600f2
f2abbd8f
dc46210f
7bfa028a
60668873
6da7eed2
9d2195f8
b4048f61
812a64d2
b30418c7
93e42a78
529c024c
328faede
cd2cd788
c7de5185
c2d4f661
cdcdf427
eb567758
d273f829
0c0f2c7a
a6593832
d99b0b6c
c79d060f
c27c02c9
96317020
eb3c2ace
55b7fd57
0bd39463
3a933a24
091a2159
e0e02419
ee7b349e
a56e6f54
245a94fd
4e4478ba
75e4d1fc
cc333b79
6f5361ac
6c45c516
39481218
758d8fdf
499068f6
eee603e2
8c1314d5
287dc696
d6e338ce
c09371bc
aa1d00ff
24746893
83c07083
ff04debf
60eb0d00
d1e2da86
29421721
e8042e3d
a4cfc0d9
ce180632
7eade2fb
8014dac6
5a6d2748
6e60949d
f501a531
388af31e
1faf09a3
2e7d3639
3b2d39ea
a258b11c
d90d2a09
7b91f054
6bfbb7d5
b44b5b8b
2b03d5be
4406d8c4
fdd96274
ee3b7602
07530a0f
b73c6b6b
ef82ddac
fbf9e685
a3721b81
fc30459e
ae883074
9c59041e
7aa49176
02093e90
33903859
a38917b6
e6e13403
d399b301
bc0dc9a6
75c03227
cb39204d
e71ce6b6
3822c718
3f5fcdf3
8e479e51
2992567b
61f64a5f
eec08cf2
2e0ca3b2
8d871bfc
3e9cb221
98410df2
c9d57c9d
ade20dc9
51393ccb
3cb2b515
d4777e28
a3fa8c71
fac770c6
db76e080
58b84e63
12f1e8d3
87fbf22a
e9def0db
a705686b
cd763150
e7a6936b
79c41dd2
a85328e1
321cde2f
30c25268
8bdaf137
a17e52ae
c4f0b63c
2259a85b
533010ca
11700275
2232ea11
49ae9061
9502711b
96d508f5
54c0e83b
5491589f
85c22560
cc0fb72d
96771c52
8a3baa1c
fb7cdc26
4682598e
eaeb63a9
3fdd9f7b
ddcf0af7
b76a05e2
f48e1bc3
59d500ff
bb2318e4
3811551f
c6ecdb91
00ff9e70
3d38e077
4832b2f5
b17e3c07
c74e5959
29dbb6c6
1fc7a760
704b6dc4
55245bd2
6219b6e9
a78b683c
121444db
bfe17ea3
a9f043d1
bf9dc249
664734d3
fa0f060e
ab8b7754
9c8d3e6e
ab60a36f
6ad50af6
81931cae
48565b9e
fcc25997
f41df04f
770014ce
d4a1fad4
5c6a2f13
d70a0cb2
b6b2346d
596a7429
e26c4eb1
bce2a409
a5176714
4cafc52d
b3329eb5
86a11441
9f53a3e1
b91e52b4
9de82afb
4cad1951
6c5c3a9d
71c2f561
c373a2c9
a26819f7
151750da
bfe124b9
7aa154d3
bae4f27b
80cb449d
fbecbffa
34787bae
ede20fcf
8bf813d0
a300526d
b46322fe
7dc7884f
d89e2a0e
fe2e3f8e
22aafa55
bbfb050d
d56967f6
a874dfc3
7af8d6d2
c3c2259a
af208e75
983ce408
39cc4f6c
a78a42d1
268d0296
0d80b89c
11732f31
c16b80f6
d7c7bcc1
f17415fe
2992004b
3992a351
10181dd9
822057ca
a51a0c0f
f9bf6778
65384bd0
dbf4d2be
ca1cbf5d
2754fe83
690dadeb
72e7e423
55953f72
f83f74ed
26f1dfb2
5701f063
18f3d3f9
545d41e5
5190517a
ec63f529
b9c68b26
6734a15e
4072a789
d60c6b0e
6aa9dc6a
c4178c1f
eafd647d
2449bdd0
f85872a5
649dbe56
9a5b6d00
49a097f2
68d4097e
2c933dcc
24357552
a5da8583
60092e39
bd8a0a07
fa5dd383
809cb294
4a8d0fbb
d4643465
74ad57d7
75c792c2
53330529
cb331f06
089a2485
e1b81ff7
49fb8db2
b4bee334
feadaffb
5646da02
2f850af5
5ad78dfa
8f9da499
a6c00966
4e668db6
a011ba01
eee4540a
c19a4df7
1a187520
d43e44b1
2a9fa200
e87cef5b
be7a1b8f
01ed67da
55e15398
dd01c46e
f6a4daee
fdb67466
e5447284
426461cc
06546e5c
1a876f19
d77a4a67
a3ca9bea
98133acc
da0fe3e8
b4dbe50d
391eecca
20eb8c6f
8772165c
fbf9190d
bcd64727
4703458e
0742ce24
b0f1dcfb
287c4ee6
b22ede9f
6741885d
2e303afc
f4f82e49
4012a4c4
03698008
3432a191
1ecf9d6d
ededeaee
e21ccba3
7c823bf9
bca3c0c3
a97c96dc
5b2129c3
5c9d7ff4
da6dd522
94a64ec8
fb962728
7d3800d6
13fae214
4660d36b
6b326405
6c24f27c
2046c33e
41923406
b548af25
6e33f1c8
fb49d041
3c3e70c3
b86b4a2b
448c0489
856637b1
1bb10db9
f55d1e77
cc4c4c9a
4f959fe0
af18b6f9
2e23197f
49632b18
a7578fd5
adf3f3c4
d980bc04
3b1caec1
91752321
e1e5ed79
e9211ac4
638558b7
99c54c5d
17c183d4
f406968f
2143ca92
d9d4a72a
1a40e2d3
e0c8e394
88fed6f8
41e3afda
e1b1bf8f
4f11e4c0
c2a45e8a
e9e216ba
5dac9505
4d18094e
90629100
e31c2502
07c071f5
5ce17024
5bdd563c
8b7bf5a6
f4a39465
a3827af8
6d77b17f
8072c722
928c02e0
eb3e2e3b
f557e528
b5bc777b
5344d758
39bc33c9
b9446424
32939f2b
6cdb880d
11e9bd62
bb412fdf
f6dc86b5
6d49f2f7
84028202
18ed3592
041070b6
41f19de3
805999b8
c3cc3e6a
b63ece0e
d2cfcd1b
5745d807
e5b1e13a
549b56f5
c74e4e20
5ec7af5a
8fb8bce2
ea8f8454
fc81e127
c34535e9
1e6b90f3
a19bf311
c71f57bf
c1ce14ea
1c63f635
83157e32
f0186141
5ba7ef14
dbb96c9c
7d87c203
b2dc2340
f1ad4c59
e229827a
fb039923
92fd69fb
ca075519
9f38be31
e12f4ae5
240ed0d2
d89edeb8
7d79a027
e0c32d75
7fd2aa4b
ca66bfa8
03000804
a8ad7000
aeb1ac36
d808ad00
a8cba9f2
0c703d0a
ec0b6b1a
b54d5429
52ab856e
981b45fc
dc42981e
8a2f3429
28ee0b65
4b0b2cc9
48530375
2d4a6d39
753a0f4f
b2a9da01
e368971c
b48fdacf
4ed6e296
9a9868b5
458b1f15
6c8cac1f
d1fbc026
7ccd63f0
e99019aa
fd6ae51f
34c7f162
1d8a146f
53474624
826164b8
fc1acca7
8ebeeec5
deab0fdd
14f1edf4
de4f4684
cf68c889
d6f808c5
e74145de
4297b616
9e32580e
d3671f81
551c932c
cd66fe9f
2f2b3c39
b7b38b4d
c6e13f81
1000ff07
50616b0d
2e793283
009c52b5
b25461ea
52355783
79bca4d5
dd9a31de
a78cedd3
dd63a94a
b075d559
777b2815
66c171db
b2353693
6f50dcea
54a491a8
b1450ab6
7b1854a9
d39d7dbf
6917d21a
26314b13
d9495e9e
561b1e23
38fb488b
6728c6c8
59509ddd
f80ebedb
91e23f35
374960c9
e38007f7
23757b2f
21f07273
1df4cec8
e05518a7
7d63ba3e
c82b4b33
ac3996db
d50c80ea
b343a208
7a8f5b4d
df709b47
3d5a31a4
6b297fa0
69a776cf
aeb77b68
8070a47d
41d13b55
c4b4cfdd
cdf966f6
ec39eb2a
1c34958f
38586729
c180278f
1d3e6afa
3ec3cd29
93176de8
63b3f514
a310cc2d
85c2013f
46dfefb9
6385ea5e
7a8c9cbc
95df7159
84aa9f2d
976c4563
24f22090
9d3f209f
fac7b676
9d7cb063
eea1fec8
835582fb
9834a00e
53e53a3f
788b87c1
e6a21572
32deda4e
93f159cc
89c59293
7e00ff24
8f479215
0752631a
efb11c8b
d2abfa38
39670008
f6e30fd8
23c728ec
8a341883
07fc641a
cc9fa309
e82bd44f
a7fbd7f6
b1748d6f
54be7169
c88d2d9d
abbb1dcf
4a0c62a8
c7d47064
3d2377b9
48afe9e3
5a09f578
03eac0cc
eda4463a
30209b9d
44df83e1
64a125fd
27218d5b
1c14d276
2407666a
353437fc
23cbf613
6364feaa
211d6452
e6c91878
ed4de331
4500ac6f
c06e340f
10ca90ac
0058ac46
c0b95112
079bc1d4
47a7c180
7bfaeb13
be8b5b30
4ad86db4
65dbd3ca
f614a634
0d753a78
8e9d835b
ab8a0477
9f9e75a9
bb4863d4
609cde6b
ebf0a751
2bb18718
06abba9c
c781c02c
7a29c689
65ee18de
37669cb6
cf45d6d9
e371191e
9f35bec9
eda8f4ac
00ff8d20
2866ae12
9660a2b0
ef2c0181
a5c79583
f2963b40
c11aa8a1
fd4878a6
c14f05b2
f21696fa
76f71694
a88b5da1
843ebc94
7566485f
931b88f9
8b3bd6c4
a34e8776
af00a793
5bcd73ca
59e57083
1fda41fb
de7e1a05
8daf605f
c984b2c3
76062cdf
00fbf304
5baaf4a9
e8c10895
77d23086
7a8c2551
a4711b22
bc1d3ebd
4263fce9
a4fa9a0a
986eabc3
7ac1cb13
51a1aeba
e8ef7fcb
e991b6a7
76a4f255
77bdbad9
fc91bee4
00dd9e68
c0708502
da32e048
3f795412
377c7c67
7445b2ae
2abec217
a1137ac7
e85613db
2dbd6d5c
11d99a8c
6be305ac
1f185313
b710a580
ef0bdf0a
634146e1
8f566458
b6db9cc2
24ed86c2
b5add6a7
afb86457
6a07b325
9d6b3f89
e953371c
f5bfe817
9c92b62c
5a9fe87d
8f84e613
9cb0d4f2
7abc0729
942ef56a
597b19d9
e34ebaa3
cd63c311
44d7a819
2c4157db
b800ff16
6e0d863b
7d7954ba
1b56d375
b41da99e
01419ebd
eaa3af77
e0784a70
3f39d7f9
f22f7688
1cae412f
db484257
aef80a83
e0a515ae
aec7587d
a1fec178
0cc9d4f5
0aa22c81
880a87dc
f4ae8862
a5fad04f
6c45f3dc
d1cf6549
4c26df51
b58b0c71
fc3321e6
e401b94c
3eea5b11
bf7b1115
879b9ba9
6a46fa4c
2257eb4d
f0e4ccda
6750e14f
3cd7bb5a
d2249e8d
e0c0128f
0420d93c
d43267a9
a26ad9ce
2aae8279
c4e225b9
64342bec
f9b626cb
95a1a46a
b91f724a
174bbb6d
cbe782db
acda9f14
eb2caa7e
1d6c8911
7c38dd76
4bdb5728
feefc8a1
78f04635
d33e7747
ba993df2
5a6f29ee
f0e44020
02f2490a
52d8a899
361d728f
465a1e53
d400897c
19e99038
dc97b8fb
9325196c
b01ad539
23fd1dcf
088d00ff
bc800248
e599bff1
60e65e45
10d8341a
03f198aa
20cd4273
b7bb10f5
70c8cb33
f0d7d6ae
fcba970f
642ff8cb
70cc8fba
3fea7f54
f600bbc2
0f741fb8
a83a7fa0
a35d8364
e01bc09d
1be98f0c
cd31fa9e
91fd6480
99c34c7d
e9475fe1
c6297c27
e7426ebc
4b65573b
570e08ea
882be027
03bdd951
e3818c2d
c7b1c95e
cfa4df06
d2857108
7286fae4
9f3e7919
b20fcc11
10f4dfb6
f10649c4
c40896be
9da8c12b
7378c0b7
8ee5b8b2
00466a07
5e99ac0a
23355723
78e4f97d
7a89428e
31225377
4c52cc0d
847cabb1
2593a102
db3df081
14bc621e
0f4e8308
af35b405
48535d8b
2ee24cf2
a18371cd
997602f2
0c07d2c9
7b86550e
e923d4de
aa5223d2
62b178bc
3495277e
1d4512ea
4ba488b4
c346bb1c
fa462840
7000ffa4
1b180936
fa480f35
c306dc8e
9369d2f9
a407bf06
e7d20fc6
99cf7b86
ab0d00ff
db65945d
8644b126
1b0ba246
a4768170
c684b0be
9594b565
9c858d9e
d5351721
1e63dff5
65dfdd95
9eb8c61f
c1552bf2
941e9b3a
5c3e311f
490babaa
a6ede66e
54c0bbdb
87d5fc51
c13fdbdd
6b83fd18
510c6dd1
f64f3c86
56883e4d
31d2756b
a7a2d88a
7912b552
4a48db74
37dee140
2bd2ab1c
8a56e395
62acce46
57f98daf
5ecb5704
c742d87a
d213df6a
5b314e98
4e917ce2
6e89f092
cdc1646d
5090b23e
758a0fc4
69553565
44de7275
d71b4986
8cc822b3
0a2c3d8c
1a0c93b7
0de403cf
f1704beb
0e15adde
cfbf2012
5bc662bd
1ca8cb7b
92a578b0
d886df33
662845fc
54ef83b8
b142fb87
5b553ffc
a85b0080
e3f46783
a4d1b7f4
aca85cd0
42a7052a
04ebea88
e3b52029
120f4fad
3f3da676
0e5823dd
b6c54569
5b61b573
ed34ce02
220830bd
827568b4
e866ae22
875bb7f0
6bac605c
f2d9cec5
d86a7fa2
393237ac
7da727dc
5ea539fe
14fd2ec2
2a5d0042
9dcf7646
d6ebbb69
4486ddde
cfef0bd6
729d7f72
286e5496
e9ea7446
f494a482
aef77b7f
1bc65408
6ac61803
33bebc19
cf7646c8
2feed51a
eed5cf70
73218959
63a4eeb0
353e702c
91be8d65
2bb5c42a
70424809
93a0571f
05bc0839
612a2377
e7e38017
c9169655
a21ff381
1a524da8
151a26a0
00d9ff3f
e0ffd8ff
464a1000
01004649
c0030002
0000bf03
1100feff
6376614c
312e3835
312e3932
ff003030
004300db
15121208
18181512
18181818
1e1d1b1d
1d1d1e1e
1e1e1d1d
2020201e
20262626
1e1e2020
24242020
2a292626
26272729
2d2a2a27
36362d2d
3f3f3333
5d4d4d41
8f00c4ff
03020000
01010101
00000000
00000000
07050600
01020403
00010800
01010103
00000001
00000000
03000000
05010402
00100600
04020301
03050603
03020005
01000001
03110200
41123121
51617104
13328191
a1c10522
f1b1d1f0
e1624252
33149223
24734372
01011134
02020200
00030202
00000103
01000000
31211102
61120341
51138132
c1917142
00c0ff22
f0000811
01034001
11020022
00110300
0c00daff
02000103
00110311
a701003f
30d447e2
46172c41
3f5f30f4
7123e893
8b745f08
21e8be50
5a3501c3
b52eae02
c7535935
2e34b4d0
88a18656
516904bc
8dc94e9e
dfb3fed5
310ac987
481d88b9
dcd7a81d
a03145cc
f802b103
05563c32
39b0b152
a1adb1a2
67bd9b5f
4a8f5617
554fb5c6
ceea18db
05baa681
a71a36c5
113c7fa3
ca600813
fbf7e3de
a56f85a6
33479449
f34cf78f
8d360092
a5b8fd3a
f5b8396c
99e275fb
9fcbd337
482b6054
a7e970e8
7ac0547f
a3434b71
73af3a0c
c07f6191
1021f5e3
c7f69c23
58b1ebeb
a913ee1c
6d28b1c7
9daec7b1
857e688b
6af45012
cfe701d2
3fcdace0
c28ad303
3ab3dc2f
8e1990a9
a8fef8a7
f2470f9b
a0cbea63
2da538e8
ff3d4938
67b45000
1768b24f
23495bef
a94dce72
a1c077f0
5fca623a
d702d7ce
07b14180
addb4008
163c68b3
e8801d78
5e947d7a
fdd47fdc
fe65f5ae
c181e86f
46b56e09
09581784
33b74027
6dce43da
1fb7b2c3
c423be2d
4b9814e8
88646755
f5ed698f
5232d5f7
1fe7fe6c
f033470b
dbc3b653
147dece8
07579b07
e10d76d6
f5e91df6
0cac212a
9046d1a6
ef09a2d1
654cf1c4
005819ac
951ca70b
5dc6a6ad
4a6ab7de
b9a5ece5
a2b9e963
447b0b1c
5b71972c
4788ca01
8dd4bae2
fe61af2a
0c7b730e
dc38c52c
8e5a3dbf
ed71cffd
23514971
1a2dad5c
36251aae
6ad545a1
6b4b3000
6dc7ee61
2338e798
2a78b6c6
680cd3e9
80404d68
b765b9b9
15404d42
01bd513c
144f0f64
a6004379
8b324cc9
08de5d21
de6da1a8
9a406309
aa5101ad
11a82abc
42d5d062
280ea9bd
667efaf6
73e890e6
edd3ad7f
9e3873fb
ffb477a9
f420fd00
3cc9cf63
70e200dc
53effafa
463bdb5e
800b69ce
09cdba13
ad8d4620
942d7760
f9809bd9
d7cc98aa
98ea7438
ac3e1cc8
00728db5
15eaa3b5
a75bfa82
7d132b5e
83865d46
cd6fcdef
8829a6fa
9c8e1176
f8f82db9
7a8c148c
b0553f6e
3eec6e3a
1b8ae6b1
1e367178
b460f591
1fb60036
348bf53e
f8d04b8e
d2a2cfe7
57ec6698
f5ed8fb4
f89a4d82
0ebd68f7
8b293f3c
924ca2a3
d12ae149
56a2dbc8
bed51c1f
22fa6164
38cf6842
c93cab6a
dde0834a
19e7d076
87536f16
2efb44d7
155ccd9b
c89867ce
3a2d867d
f24a0cf7
d12e309d
3fe2fe98
2bcf4403
2b19775b
517ad9db
1e59934a
e3ea605b
bc653fe2
f537ad35
cca7921f
f4022b3a
e91cab84
01bc605f
2dd5dd23
8f1337f4
a29fee0f
d90cbec9
36983850
81fbf759
f3596943
13473785
3828f361
5a392c55
393df67f
bbef3304
a8540aa7
eed68fcf
643bc203
cb6797a5
9507221d
ae4c588d
e84735d8
0037b626
0fa58da4
258eb92d
fef6ec0d
293a8163
a2e4a315
8459f8ce
5a8db9f2
2ad5cb17
5d4c7b84
05c1511d
9a23c453
a3e42038
630871c3
432a8277
c212bc1b
e02a7580
a09538a8
022be82a
a1952abc
cedec721
7faad5dc
44c89ff5
af0f86db
10dcd3ae
2e3fb49f
d7de0fe4
52f0e337
49fa6625
81fafaef
d9655280
2a8faa77
fafa9953
dfa021f8
a2fcf055
9cd93917
aecf0e23
a40ba95d
8d982813
ff5a735a
a2e9aa00
cc827b6e
bcca4dd0
346244bb
62da2e17
c162b9e7
7f6e3977
ce33ac45
e877ea1b
c4c99db3
bf38c730
7f6a5472
7cc08023
ae524d4a
9d1e74ae
d10ae411
754dfd37
6dd1d3ae
e0b44a75
5c5bb79b
6646d573
69c103b3
36dd8b71
98a3ee7e
2af7873e
7cd386b9
48afccc7
ec0957c6
9c77353f
9ec38a07
7322aa1d
c8bc44ea
f38e481a
5d4b17f0
c459a45a
fe26395e
f997fd39
b753933e
2e93602d
57f6da18
01a8a0b2
0436ab67
9eeda16a
fee9bede
7d80e692
1f2dfe6f
7699a2df
904a615b
9fec326d
3bf1a1ca
815e00ff
ff312907
b6cc9300
4660ca6c
6ebf536f
854f8983
83dd8c38
c61af305
bbded137
ae2d9a94
72583ac9
99abb55e
6d204a57
47562b00
92046355
3d50ea00
4502787f
3bf5cf26
ade93ee0
3e5a9291
99b451a9
29aafe98
67066fdc
631c277f
b5243af1
27f71537
0beee2d4
e764df6e
45877599
2b7dcb35
be891fc7
ecae8fc9
6dd386cf
24ca82ce
fdcf3df7
07b5aa7b
ffb37286
7dd85600
00ff7ed1
3b2918dd
fac0b76d
1a08fd5e
45a58e37
8970aaa4
31aebbb2
981b9329
0d261680
d1b76f51
00c7eccc
268b6e89
7a7b86ee
3530557e
0544eb29
b5950443
e5a02b73
2c5cba78
144f0978
04044773
dfe651cc
78940c04
bc3b4333
dd184a11
1eb152e0
16d04a9c
85578973
b86a0565
43cd552a
860abd39
623c4695
f7a602d7
0b8fc4c3
1fa48384
072aeeae
adf64d0a
d431aac3
6789f20d
106277c4
fe259b32
ca532bcb
cbb7814b
140a0d8f
8a4eb73e
2db3dd41
c1c44037
1f953a9d
18b6c1bd
5e119b68
fa61d139
c85cf02a
f5a87a6f
ab18d9fc
7c548fa4
99b52ad6
8308de94
5ac38a07
e1195bb6
c721f936
4730ec10
96811dc7
baad6a5a
b7f4982f
a1ba90f2
d5755838
5712f754
77a0c14f
24095df1
7db5ed73
60a71e23
bd69653e
a3956357
acd2fde7
2d3a80c0
a86f896c
6282e144
48ba3cb6
4793271d
d3ce295e
63d3e761
4ed612aa
88377562
7501ac03
5d9bdac6
f330792d
01034927
1a9b4ac1
c1e7102d
8d6ee981
5cc2771a
6302a7ee
d78ed937
16343268
2c3ca4e4
a9bb1aeb
004ccf4e
16829a56
d0a2d24c
b042b3eb
bab55819
271801d4
24604663
f7b92594
445bb256
9f188e79
ede93ee2
419a794a
4651f5bc
c84b9ee1
be7b2c3f
e21bddcb
2ad5eadc
cdee3938
a007e9a8
de6638c1
de6fae93
39f11884
e9b41b67
2a3d51f4
74d9a4cd
ccaae998
f698e0e6
30206d20
a26ba001
dccbbd8f
771b9ac1
417d707a
9737b9fc
7f7fa85e
3f7775ee
e9f86fe3
e235e28f
7b614275
a1b95e0f
8bf89e65
97ae5549
695512ad
86d9da9a
4c6b4ba9
a806a653
3b4f691b
041449e5
3b9382bb
d91f4ee1
5a015bcb
d4285ebb
952b5caa
2d47cd6b
becd23c4
a3980908
5908bedd
d6500e0d
908902eb
8602efd6
2b7174d4
4a1c5448
ba6015d2
b4563557
8821c4b2
b48f11d0
d97437bc
ef2d4dfe
645c5242
1c532b99
9be6e058
43882383
9e07b76e
0a8758ed
9abba463
829f098f
6dd6df25
71a3b677
d1610673
910dc5c2
ea2c6c95
7219cc29
71c57d52
f404c194
346bee54
13b2015a
1ed7dd7b
0cbb4298
f36cca37
2a350dd7
b84ec2b9
0571cd25
7a1a6e74
c5518508
fb9c265f
d6e9bc76
ec708a56
3cc83ccc
25623116
1e1a156f
746c10c7
e3e9a6b5
0303080b
b065c328
e1a88073
66e37f77
2e79e6ae
6a10bbf6
034bbc17
39c70dbd
bb4bb9d3
5da6617a
1df238e2
fc3c8f02
308cda4f
8c447ff3
a5250ada
0713a7de
c14107a0
b937301c
d6d0ac62
a4851ac8
f19d32b8
d84f3c2b
9524cf8c
901e70e9
0216fe64
b15770f2
66b187b0
84db7426
2c8b34dd
24424cac
c8e55325
52ba6751
0299ca20
725af702
c329b3c2
a6a0bc71
0c1d093e
a3c2288e
78eefcbf
1228bfbd
a2a4a2b7
d63e47ea
0f7e7aa3
73c09fea
245d00bd
115fd095
0a38d275
80d1d2ca
940bb3ea
cc4f6fef
2b8b06a8
2ca54dc3
8b52e794
6381dc58
d181cba4
b7cc853a
7c9a7c75
4e95ba1c
8d15c455
d92c5c69
f33aeb8a
84b8fdc8
00c1b779
ed1fdd34
281908b0
776f8887
73a84481
6a438175
b4223e39
8af89c05
2c4115d2
b750b557
8eeaa6d2
fa49d0ca
09ac43ba
a450b283
13f58eda
4704d29b
e8847649
92bf8db7
22127ce8
aaf84947
1c398a2b
3616032a
6f244430
61bd6d82
1a0319b8
bb9c33c3
63c54fb6
cbb455af
e9e52081
4a727870
41a3d7aa
2169cae7
92cb4ffa
f5792f51
f1a34643
df70ec2a
d77347d4
49aa62dd
f9717112
97414505
8a9ffe28
a37317d5
58744c00
d4d1cc49
74e9624f
d121d7e7
5255bf80
0bfec2b7
882f32a7
2ce61538
26f7148f
f41f7afb
a7e40cbe
41073de2
335bc9cd
930b86b8
2653efe1
302968c3
dfb4160b
9a7deafa
4e2dcfa7
3b8e513b
72edda32
9f60d98c
7e637f0b
15cb3ae5
a6984603
5c5a198c
dd124a6e
04b3996f
76577508
d0e79937
b153e428
29b3e20e
1a9cdc0b
dc2f4131
c85c92d6
35d0051d
8939714f
d5eb3127
67fdcd54
74616517
9ae3058c
0bbeb22e
40ca332e
4ca4bea7
95a5c83a
202df118
769d62a8
94f130d5
e21faaa2
81572836
8f3529e7
6aa1334c
6a53cc2f
5c9814cf
a50900e2
73fe8665
4140725b
22fdfd3b
541034d7
26f7bb7b
7709c4bd
db1d0de1
d3903e81
6f7511d2
61257780
d8b938dc
396f8f22
69bd519b
53a914ca
dff6243a
47581d11
85fc13cd
c4f3203f
65593a12
719d0936
5be93deb
ae024fb1
c2d61198
1ce4029c
b7a314cd
1d8d95a7
61a33350
20a23e39
56b9554f
a0b2172c
c557ee58
c75abc56
558b2a04
c45ac9cb
5210cf62
a300d746
52509f26
21d8d45e
211134e6
44b1d8bd
81757be8
e4463c40
17be8a7a
8056c4c7
213123a9
364f98b8
84daaa2f
480b86b1
9f8813be
5479b3ec
bac77c9e
0b0701e0
d5547158
0a3896de
2de40863
c9d37dc8
69d7adb0
b616ad1e
7bd4dc81
7141ea69
4ff48f39
c650f0a8
5c5e7ce7
dae5b2d6
cb421af4
dc54ddb9
e037e73e
050b800e
972c1dcb
e1fe4c13
9ac7e9a8
9d540fb3
4bd9cba4
f3bfd34c
cde174ea
39224156
ca6b1ecf
56669eb1
0cccfa96
0fea4066
ae926e45
fc91d3a8
aa68a4b2
02b34366
1613c362
c43f0d01
4f34e070
35c7f14a
825c09f9
98700546
f59aa8ed
b8187003
3b1403f4
b3c8d974
79ef36db
7466e06b
fdd57086
859a29da
0300343b
f87d205a
4a658794
80c0b604
1f8c8ed6
ba79d374
6d79461b
ff70d420
fcd45100
2b7f3717
5c6be8ba
d8cd7b47
ef3232a2
79e6f58f
ad290af4
745975b7
29f33893
4d463dcb
4ef5c4c9
4b704e1b
e1318dbd
9869371b
757a0240
f643eafe
4ba2999d
ca6560de
ea4c221b
b1a22ded
58d169db
1203b1dd
5466d13b
bfc3089f
733552db
eb68a0b1
618ed063
a2206829
4a0402f7
19085948
b14b9028
8705776e
14efa5de
77a0b5a4
e6eddb4a
ef290e2a
939753b8
3f63a338
cb2f0bf9
6c6983f4
a6b767aa
0388496c
f7a9ea58
11cfb506
adc2a8a6
eeb90932
60d45d28
e4f25bf5
2ea0862b
dd1e4608
5a1dcc6a
eadbfb50
56764fed
3d8233dc
e5e489bb
73d8709b
683e12f9
dda25c78
fd55cbf8
5c300cc5
2d3a4df2
4f69e7ec
5aa55035
5610fc42
472e96c1
4335c4b4
8457dd9d
2f5e68d4
5f71ca97
95cb172f
992a3caf
8ec6145d
2f38d5dd
a6214f6f
b49d14e2
86ad28c0
4c5b4ae1
c466f602
58f78752
dc21f114
c4c254e0
6e457c7e
7eb26e69
f78c084b
0d0d6fc1
8fe11ef1
04bd0a6e
d386fbe5
e9a4b1f0
d62a8632
80c1e6aa
02d00027
f792f76a
18ada135
9f9f1b97
f6ac27c1
937ec3b7
ba003ff9
ca21fd38
1d41b4b1
54b4605d
118f4073
754b0317
8b0bc358
b9493049
b4c09ef9
b88b65d7
0f26883b
d4ba15ce
4922b249
54d65632
c318c0fd
b5c29a4f
c39da7d2
742bf40e
57d8ecf4
005a8339
ce5f3ccc
ddbd920e
0b1a6b51
8a7e0b44
427d54da
c3491bfe
ae2792b7
a57050d6
a34e1f52
878e7966
e7920a4d
e23157cc
7b2705a3
8686d46e
3c97eae0
a0f8349a
5611adcd
095a5cb6
4800ff24
64c3a9fb
ac8fb1c6
13636bf8
7bc56880
4bac77d9
5debd684
853dcd7d
f049e40c
74ee6fd3
2caa067e
71d6476d
c6b9cc7b
fbb75849
2df7fbdf
b64d9170
6ba43fa6
b457e2c4
839ab250
26767761
322551a6
c6531886
24a23315
b2c20b11
e4d2ca35
f4c8f450
476debad
a1746f24
ccec9ed3
7feb0854
a3504ffc
41bdb35d
5eaf7b49
0ae98fd9
9f1a3f9c
f546f13e
10781f82
66a8fa53
e3d3b2bb
414f3e28
d314f18e
34c56d6d
2531a791
bb62a434
73aa300f
fb9bfee7
dd417d9b
0ca5fe6d
afd17c34
cf6936b9
e5507e47
d1a86706
e1bb65f5
db3c72b6
84c6ca53
6f52b050
9c2b31c9
74e55aad
95f35ab9
d658f9ca
f3021097
3e7abbcd
6623b963
a64230b4
a14d318d
73250d6e
cf74cbf2
a01e6dca
84a74da5
658bea28
71bb49c1
6f862e00
ee917c62
49d029b0
281558b7
73431db1
5dc13d19
6e2cb89b
adad15f1
fa9c0ecc
3223032b
eaa71ee7
7cce2716
03985ca0
a433eb9a
b3d006f5
a35e1a97
a43f9c77
e2eaca7d
7fb2e4e5
04a01bc8
6b2bc677
139d9e9b
94679ad4
58baf3e1
8c1c09d2
329de2f6
040e4b0b
4c9b0766
054115fe
458d9932
83be258f
b3c3d798
24823711
aa56828e
e3aac894
8adbafa3
9b4e77bb
96314d8b
214e37c3
163a6f49
2b66364e
e3df4583
03e2d0ca
1dfd2289
04392613
a88efa30
11003966
f7bb1d15
d95c6e0d
22f9d741
b7a5b213
bc847b68
fe4847f8
f8a95a5f
e5ea63c7
b6b76da3
04319db6
3b331087
04f63819
4d37dd9b
f3f92f65
0b0436e6
f8c0ad01
4777d5a6
5dccb669
a4082a35
bc1a70d0
12953afc
92b897b8
3dc9b864
df8c5b49
85afec35
446cbcd4
d443f194
44f1f6ec
cc25f16d
38351ef8
d5d44662
c3e84285
4b895680
67c25ac1
0513eb8a
c818352b
88e271cc
4656d09c
79ac04d0
8746958e
bf22055b
27d30e70
6c26125c
b19eda18
5da89f36
20a600ee
eef80808
d7650b6c
942a86fd
83abbf0b
3545d007
e82419de
e5516114
a23a2eee
7feae6fa
6b9a5a66
384cb6a4
629a8a1e
9ee2cadd
21e904f6
0e75406e
24b1072d
e272eaf6
0ebb894e
f40fab7d
664b7e90
7d4a9eca
a2ae7cea
21ca6e9d
5fac8060
3b40b968
7cf1e2e5
ee29c7bc
4a679ece
6d368d44
75e72086
83097b0c
35b60a1b
3c63536c
0f2fcba5
413c34c9
027c9b49
a462a88d
5f01becd
424ecc92
94f0ba4f
728b04f8
91301524
f85c9019
8875510b
f74f0018
6c70545e
c427b7b5
e692037e
96e9f2a1
b2af1ef5
340878b2
3162061e
3312ea03
d2a86fcd
b3320f1a
e124b2b5
8ed6253f
4bd05a55
da9aeb67
711038d7
e5a8d32d
326b6cc1
f345b36d
aa6ab03b
11e33a00
2e8a877e
d7c26c8a
94cd807a
98b4417a
762ffb88
2d57479b
986c0135
bd8e836c
6a1a2bcb
70ca08b8
b5c7a881
e650bb48
976890be
8136ce5a
d98bca8c
e1f9ae75
fa7b1366
fed76630
e1a86636
eb061b94
522875c0
be345fad
9a315bbd
6facfd75
9728f733
a8bcf376
5369fa72
fdcce99b
ddbd5194
3ac5abb6
e1a9f87f
e7d56efd
4f02c9e1
6b88d795
03eb3e75
51713beb
b0741ef5
408301d0
fc4616e8
aede0155
49556be5
389c859a
841bf084
99d2e284
5120dc34
a6b412f1
165b290d
8c4e54b0
e7730535
b45409b7
b42875ac
db3416de
d6421dce
9036cdcd
29269449
e5a97eb4
dcdcbe3d
8c4471cf
a2709f18
1a41e661
50dc8e48
ca78e7c6
79c565a4
32d89e52
666e4e03
da42ed50
11e82e2d
36a8feae
d5df1f48
9e9b9ac1
63055408
b8bc6ade
ba60acea
738c4fb6
995df92d
74b15bb4
8e04d3e5
251e7525
affde228
c81c6dab
4c5714f9
db5f0840
ea0fc7ae
3e051905
a5c7a97d
e5da858b
cb57ce23
cff3e2c5
6fb48b94
62e828a0
6cb5b314
9bf32930
94ba2dd4
ba7a21ca
9ed3ad5e
b64593fc
1cdb430a
c8407f14
6e00ff08
88af9389
d61d529a
77493a05
c4031458
ba55db72
36ce5959
e4986eea
8272de73
0334e662
9dab8254
938e049a
0c5d71d2
bc722927
987d5731
2a3fdadf
41232299
6aafb83d
70e87189
77bfc959
9f6374e1
e5cb0f47
1b6ecad1
24698e9b
152cdb1e
06418029
e9081200
77a0a2a2
9cb4c796
aa56d81b
0b04916f
dba9607d
e642c51a
73fa45cb
3da3789c
f7cafc8b
041f6673
c1e7639d
69ad310a
0de210b4
7fbb10b1
9da3469d
06ce5e4c
1f79b225
7216359f
873756ed
00beed5e
8244cd7f
eaf6e6df
148d687f
bc5d316c
2e0bc3c9
c6ad2498
df02717c
5d354e96
457a0503
f34eaadc
65468b7e
105ea581
9596386c
4a079a50
46ac3907
c73a9529
2aae295b
d56accb1
b20f25b2
58d94eb8
4a953e15
7f9551b4
2979b1fc
16022a8b
e913f082
416e0ea4
6f1fd56e
682e662b
d13bb0c1
c2987af5
497eaa8a
ca091f25
91e1653f
67c1adb8
6ac52fa6
c391ac0a
ba5a7826
df58c1eb
5fdf570b
67a12235
b95361b6
87506a18
f200ffb6
342f22f7
5d164202
5f6f3a8b
2a60be2c
6ac74ac9
a5aaf4b5
e21bcb6b
44d1541c
50f03645
eab9ddf6
485373b4
ef1d42b3
3b7d06f4
52252e5f
6d2180ea
29919f3e
3b49213a
340a4857
7d147273
371bc1b1
5d9a014f
0df59959
3ee0b81a
4b0813fc
47b80077
c030055b
9781fbea
b534dbc8
fc9dc3a4
3aae1eea
1ed57e34
aee62a6e
d990f470
8f6c4318
05ed8077
f2826d5a
24f4a4dc
76eb8ec9
bfaeaca8
cabe39ae
da13e862
815d3e15
6365b6ea
299f1bd8
d903f5b1
b1725a21
cc98b3a1
1c013f92
062f3a13
5bc35b9e
50c71a0e
823a65b8
ea08b6ac
a5243f08
931ac7b2
47797e94
6bcdc344
07b4bc72
3c2d801b
dc0c33ca
37d61245
f3b8dbc4
56f7aafd
96cc2171
139b6893
a4381ccc
de38dd34
d90f3d4e
b4803111
27b4676a
ee32b2bc
05a98df6
2e57c98d
d23e9a6c
8db5fa63
8b20a550
ce551d9e
69355b63
ce98e880
0259d3d1
01aa2be1
74b0a802
8fe1e8c8
8e6abf68
f89037f4
abd67fb9
e6cbd43a
ca59f1e1
d8e20d24
d6165216
cdb48409
9854442c
a27d88de
a8e9881c
988155f2
606ad131
f836b232
7d0a6d26
7c68d3aa
72716c2d
4c73025c
a3dbf642
87635186
403cada9
c73e7748
6409aeb6
ddf477d1
057eeabf
5bd63114
93ca5481
1ef78028
4bdab9d5
7fb4738b
62b45f36
a51ee010
2fa8a9fa
dcccec7f
32004a4d
35b825a6
cf6300ff
037b17b5
8e068348
8373c52b
20702d9b
c4411087
e208422a
509985dd
a0851ff3
c85695b0
b87a867f
7b83f0a7
9c0fc413
aef95ccd
c26ad909
ce2b61ea
1568e106
25cd4a81
573c95ae
18dad3ad
ac816b7b
a8fb32a5
93e8daab
94a2bb58
5dd914e2
5c8ef2d0
debc11e4
61329836
7c6edf69
d40d12a6
f7b35629
c9c6252e
d2e4d9a4
a63ceded
00c70e51
0396fb96
f0b0678a
b8b15785
a6dad20c
45103308
cd145ffa
54e0dc29
f730226a
7009956a
98a94126
d734a61e
06420629
aad3c605
0d02f727
06e4b84c
ee009dfa
173c2118
9c9c0e6f
f69e5ffb
d15560c4
cd71cc2c
5171020b
60b428b9
70304a66
044936bc
89b4e2f0
4d7d1278
b3f02730
9727511f
12e67bcd
ad2f7c2f
b2cdb096
10c591db
01a47fd1
24387273
63d8cc94
33b6dfa2
db290e54
b63c1e0e
a94fb336
72f907b3
95b5e0ba
c01ceee8
506dd260
087bf10f
92201c0f
0cf7ab38
86001835
f796b8b8
ddebd269
b536aab8
aa7ad618
20f0c692
41969e49
f39191b3
5b05973f
0f96d685
6b3e1017
372909c7
38287cc9
9890ce04
3b612258
af3cc4a2
71396302
4f706550
a2d18ce9
5bb05551
2ca43dc5
5245bda5
219a4c73
0b280b6d
4d752a40
525a4d6d
ad34b7a0
30a5e578
539a4969
05689426
1a4d693a
6a3a3194
239914a7
07d87bcf
8f69eeb0
00f94753
23ee7ed4
36194a5e
89f52bec
89b4c001
82791004
b66f31bf
a9b86de7
739bf64b
dc920f07
9da271a1
c7348aa8
724a7b22
316cd1b2
d45aa0a3
4a2ad52a
d64aaab8
52b79033
b3006b66
a60da5e2
719836cc
ca4189c4
5e73729b
4d137dfb
798a91a4
185ac050
fd9d2120
4f852d7f
c9f203d4
6c957b19
3a082def
578d0934
563d7166
66111570
7ac43d8e
f06f8f56
4dfce685
05c3ce35
ac3fb14f
3c6e956e
b859a229
0ca546c1
74544cef
8c2c945c
8e8acdb7
42891fe5
85890320
27a7c3da
c1b5dd3e
f03c17b7
66ce430b
cafc3789
05c048c8
346f30ea
d5f0f58e
ca1f0474
bcd3ade9
aa312ff7
12a7bc7c
f444d107
83cd480b
0d258e89
8c04e634
890ec745
b5522abb
a6c509dc
db1e7922
7e388da7
41cc21e7
d6022d73
b8adaae6
e60658a5
b62847a9
3596cb58
e65fca8b
60c7dc43
c5bf9f71
1450dc67
73700eda
b41a6840
10687a6a
297a9be8
a392d135
2d139920
5567c2b0
c72dec8d
597177a7
be2cfce6
f58e48ce
241ada39
1a624aa2
7e6ad292
2ad9142c
125430c2
98f684f6
7a361280
89dc13ea
b8a810da
d4a50baf
2d94902f
4b696e05
8cd5d842
5a4c6935
bd958652
44071aa5
c272ca54
f994e986
2c8a5785
ef49d48c
6df37fdb
21e381ea
3e328887
0709584a
a81551b8
c7836373
6c94f677
c04ea0ba
451710cc
c3607d61
a559e10b
2b4ba773
a4aee042
add8571d
5c42aa63
a691a938
880ab629
fb44d85a
e61cf56a
979047b1
4c80c41d
ee455432
85b8b315
925fee26
3783729f
a5c42535
38d7b3ee
eac6a5b4
ac023a87
7a9855bb
17a4aa8c
c9780f69
fb2478a4
19b85914
57081ea9
3daa2066
6ec0279d
84cfdd12
51c24cf0
2837b5bc
e15da254
02d4e390
de2a0a84
1020079c
ac5df2b4
edf3723a
749d40f4
2e00ff5d
28d8a50a
7c213dc0
4cdc553f
82868bc6
6f8c974d
209ccd41
2d9ccfeb
76b376b5
b1c160e0
0abddd6f
228bd047
95ad355a
70022eed
6cafd8d2
2ed1a7c5
81e5b824
963ce9c8
07cd5417
2a4db008
21461890
995b1bd8
93120fd5
5d2b7b4d
68622531
36298892
6c746512
b629cc66
656a5517
3a5ca911
f43958a3
a8615255
7d51ceec
d750bfd5
4f284f6d
2d30b39a
c9547b8a
c8d5eba5
a532a456
f0852b78
4a83695e
d5520ade
613ca5bd
4c7d0acb
ea9486a1
d458959b
2b2041b9
1d0409d7
b4b3da6d
855a25ad
4971f7f9
9cf6a8cc
693ee25a
906a2e41
4a96dafd
9e78f4f9
e11664f1
55350b2a
00ff5ff6
d2989a43
43e95edf
528ab0d8
72829b6c
3bedb699
eab0c896
8334f689
ab444f5e
b2ede4da
fba565e1
441a6da6
f6ae72dd
6ebaf7a5
cd508872
d58ab94a
70bbddbb
553c52f2
efa2e398
158f465c
82c56497
400572ae
db44a3ba
0000d9ff
e0ffd8ff
464a1000
01004649
c0030002
0000bf03
1100feff
6376614c
312e3835
312e3932
ff003030
004300db
39303008
42423930
42424242
514e484e
4e4e5151
51514e4e
57575751
57666666
51515757
60605757
726f6666
6669696f
78727269
90907878
a8a88a8a
f9cfcfae
7b00c4ff
03020000
01010101
00000000
00000000
07050600
01020403
00010800
01010103
00000001
00000000
03000000
05010402
00100600
03010202
06040402
00010103
00000000
03110201
51122131
04617141
22329181
a1b1d113
23f042e1
f172c152
01010111
01010101
00000001
00000000
11010000
21024131
00c0ff51
f0000811
01034001
11020022
00110300
0c00daff
02000103
00110311
5a01003f
5002d187
ebe7136f
7c811be8
902f6881
82868019
4e2c52b3
4d8ed0f8
c38b1808
92382e49
9528b8eb
00fab986
2a2c3c32
b4c60a2c
dd72665f
da516b0c
2ee14c4e
db12015e
e35b3164
8a9d1115
1824e3d6
82869106
81b03ddb
b165d91c
40d83642
986551cd
3f5dce4c
9d9f8160
2c1aa558
56fd0272
18bce63f
d37e8926
20d980d9
91d1f6a0
7c574f7d
251808df
dcd43490
37ef3dbd
48524b5e
783ca2aa
57d49565
db89ec8b
dae21816
c9bb543f
3b461ff6
e4635c52
8e6cd931
24b5929b
b59cddb5
d79aa619
cda62663
aef81102
ba26e351
89c38c36
569f94bb
e41aa1c4
da108ed2
b4627231
702f14f7
a9b422f1
d7e6d450
78830440
893ce880
0a645235
6c810ae4
6808b482
012a2f28
1714a161
c2280ea1
e8fe71ae
17bbcd3e
d99f7f7a
33b9278f
0347b351
662021b9
b2129bb5
6b62aca4
4b0ccb1a
538c7d73
88f8371b
505f36f4
b1dfb7a1
f6ac18a1
978529cd
d89e35a1
152d3ac5
21846dd9
8a55d19d
f05bedac
8bfcad1c
f6b7e49a
bfe98a3c
3c92ce98
688d1155
e99bfbbd
3c2c9b22
1e9f8d45
b64af208
4acd9443
c767f9cc
03939f1c
e09e56b9
f4c9abcf
7f773dc6
88d853f0
edb08c19
22ad0907
560ac748
b285e20d
64554445
f8a0915c
3d4295f4
a840d441
a1023187
15c818b8
28051903
d0a0b804
f2c20a56
3e0ed1a2
ffe4caf4
4d13f200
d4997e02
894453fc
2a25b125
ad1a683c
b1dd16c2
6906090b
4566a4b3
168d18f6
66478c76
76ebceb0
2ae4e767
e54cdce5
4d0887d5
b58117f7
8cc04bca
6cd82bf9
f18a36f2
e3948f36
1191bbd4
5c8bfb36
bab0519f
2fd29c9a
2137bd52
479e70ec
b2afaeb5
e3505c26
7d775a1a
f81b80df
ae4b367d
bafaa0ef
1d5a2a9f
a9675788
0d04971c
e4c8b4a0
533f0f90
8cddabfe
2a6af3c1
3779a6c8
73aec4ea
316c739f
ab36a937
27f10d93
88646f37
e6fe3c93
2fda3e49
cee61704
dd43b8b8
535a04fe
24035713
dc82c4ac
0a61b731
a1788433
d34628ea
3c39e898
e031383a
01620e22
2a00f220
20673083
15640c52
67d0f488
69052c2f
33704971
69f1c59b
bff726f4
4d722083
386df3f4
1652007c
6a0a344a
a42207c9
d0d0ed47
9c958d57
e32a0695
c3a8a414
c3385029
52ad05c8
0b21f99d
7d3a5391
be9e838e
e6a7593d
d6a8107d
5b316ebb
7b00ff1d
e6e1710e
4e2d7b93
f7d99320
5a514c25
5ad065bf
8fc73124
b247b565
b66547fc
d721b264
d4886159
122c1a3b
684ba89f
4100ffee
a28856eb
6c3c8b6b
7672726e
22148edd
7cfb04c1
45c97802
0812656e
fb887d14
07e17f3e
c0d777b7
539ecd1f
02ba6cd9
d50aa467
a84767a5
e85a33ad
20d5584a
926d1c1b
aa243544
3b2dca61
a852233c
f3acb8e0
200fca51
00f62001
d620c7a8
c81a9840
d2e8a80d
052b6950
a55971d1
31a01103
bca6eef4
498d04f6
a30db4d3
eb2d51cf
2e8147e2
d7b42969
3688bf75
09dd5469
678a3de7
cbb60924
4c6b4da4
33b9d8a4
ee4585ae
de42f37a
6adf8cd1
81851dd3
ee2d2c86
f18ee8fb
97dedee2
b04beab2
1da96b8d
582424aa
1cead5f8
5249312a
0423dd34
d8b76766
03e965c1
1ad20c17
21c45019
6716d114
5e003289
5b193ba2
84615210
09d8d09f
1d5d982d
00c3b1f1
a0e3a3b3
a3342be0
930bee30
38a6e131
a3520bd2
e6e8501c
45677d2f
5a637034
75d60c4e
e8479e67
8300803c
0faa00f8
2881bc01
511b9039
9f4173cf
25a8a4b9
dfa0e885
10f6e414
a30e06eb
eea75f1e
eec5e16f
ec342e51
5c429346
ecbca4f6
f67139c7
83514a15
8da256fa
4817bbde
f9a5588f
c0ab3d94
7598d5d5
73cf4947
33ba4565
67318fa6
cd21bc51
6a452df9
6402dfde
f08a8fc3
4fec5ffd
b10c896a
c1ebade3
deaa4374
60658b86
1fab4c96
46e89f9c
283943a4
9c4b00fe
e619a0bb
cd52a9df
2fac7427
02127fe9
4ae11ecb
1143e869
54a19692
a443903e
0b16c6d4
f8a48d45
df3063ab
6c4e4092
dc23aab1
417dd399
50fab8af
ed665850
4d771885
568e0279
d8d76012
1e7a8127
b59c5166
a4138e15
c05d611d
54304ae4
3e340a90
f4acb889
e2b36381
e058c3b3
0d8f8baa
925a3162
5a323246
74305e92
90371061
00b20727
5eee373a
52d0dc7d
98076d46
76d9939c
dd8b7133
a76599b2
7924e1b0
6df32845
3b7c7d2f
ddf2c490
6799bba4
39f5cd91
f3f66d4f
2d299f2c
acc4d32d
569a5af2
3557a9e5
8511f6b3
3d0d365e
72c62b47
79843170
6883f8ba
a71b04b3
93f8e9dd
43c01734
b0873f8a
b64f26d3
f4cf7ca9
bc83ae39
b5ec3899
50a688fc
b772dc72
d828241c
243b968d
8e8f4f3f
899fa6ef
00c50267
cd614cba
bcb4f208
622f2845
0954014a
1f662b71
a2e3bb53
7bd4e136
701a6e99
1c1bd42b
e614fa4e
4409c356
42377117
876158c0
fb005ee6
7c718f5b
69763ae8
163cd8ad
184cdae6
1ae71443
40ac12b9
7ab82bac
e3aa21b4
f1f1e141
0f8faf38
e1794d8e
30c6d049
1af23c72
8a8c9d44
3d6329d1
fe20054d
6486e041
e6fea3c2
e61e46e5
c24aadfa
6497e672
6b524a0c
bdb71af6
f2c4bc2d
62746869
33bfc61a
d5319a44
bf4ba6d1
23426ab9
264c7d6a
9e60abb8
2ebde536
e49efbfd
d8624b8a
9e007fc7
7be94769
bc6a12a9
839d0446
5fded51e
3c8e1990
184ee4a5
edc94992
c2bf1ef8
62cdb9c6
d525fb8d
93936291
6531abb7
9fa6f7cb
41eca165
0499a051
f1100691
43223a13
b66522c3
2b463614
6dc4d666
2dee3983
88bdac43
4b720fd6
2913bcc9
467c4f9c
fed807f2
20ddcc40
463d0627
91d0f990
cc8f346e
7cf39c8a
60f7dffa
97b90661
410eeed3
79b4465b
06054905
ce89a108
e8e4ac56
9c9cd7e4
6725169f
79846d9e
292ad930
8e1b698c
537ea67d
32a6925a
9ba48e3a
875ea103
a1833cc2
51514236
665dd6d6
2bada937
568f0c2c
d5d17a62
dff13db3
6375e4bf
a3775697
f0a3566b
d2d22116
4105febd
16df2805
52cdde93
2ef3535f
3bae93c8
cf142475
a5f6d29f
b06d18d4
4a73308a
8730bfae
de0a46ed
3ff889bd
4681a14d
d9c47d3e
5d7854f2
ed93a58d
f277efc2
af44faaf
d563737f
24417574
82eae841
3c3c2d34
43238443
9ce84254
b1e6051a
ae902b9e
6822d4d2
cc63a0c8
45b29271
1d00ff73
7b159608
f060cf9d
5c80c400
c914ecb2
6e3718d1
b5f6c4c2
a6dcd9c4
9080c325
843dbca7
ddb86398
6ce0056f
f5441ac5
1f168548
e33b801c
cce3c3c3
adc43d72
6b4c8388
a3c73460
36d28a04
bfb64413
4c52c724
93401b81
1c565f20
840ff289
19112653
371e35f7
97732f5b
83c0a2b2
df8ca857
239db125
5a2de5ac
037f531b
760f5562
9b52a855
5aeb7b2a
e5c6e31e
2e95b157
e322a14f
5544e3b4
fe583064
05f6b6da
29572e25
82b4bf68
3dee8f5c
8c228ab6
2f9d14b9
a8af7e95
c981990e
00ffb6cd
514446be
a4a2967b
82c75dcd
0024831e
04432578
27b2462b
92e7d444
14374629
1ab94d63
e904d2d4
1120140f
1dbd1f83
52e48941
56a8f1d0
2aaaec80
cd1f02c3
63a9c02e
22969d7c
339d39de
1de94c47
5f1c2575
6805788f
f1a3c317
98ea890c
e4ece0b0
1e9f9c47
f1791e1e
115be322
5be32cd1
1e99d213
e79a1e9d
90c424bf
0ff147e0
f0ba12e0
3ac8214c
d101cc12
4916f2cf
c4368db1
113abb12
d393622d
5af6a4c8
9e8bce99
ae517538
1d8a0686
a4067ed2
76d758ca
3bf10cb6
28b8ab96
6fe75e92
fd715b94
eba8aa88
11fe65d4
00ffbbd3
ce766c84
01f2b391
bd4707d7
bc79874a
5e0466d1
c858e204
e33e6069
159bc828
011bd568
91da31f5
4bbca53a
33c5d8fe
06d28e45
4ab28fa8
a60f74ed
8887a9c8
193722eb
a3aaa8d1
a2235a32
22f1a1c5
e10e66a1
f9832180
0a815c04
b2657cde
acec58c1
96d7a8f8
3aa2492d
b9821e22
05066922
52707c76
c8ef24d8
8d936491
1f54a391
385d0d62
5f491733
5bc09897
0786c93d
82707b4e
97f7dda5
1e91978f
0d2f574e
5fee01be
5a4bf2f1
f13a2ba2
a62ca6cd
ab9a948d
95ec96f8
38131c6a
dca2abbd
61cb27e1
83ded94a
ad53490e
fdcd30c3
5fab9634
eac9bdc0
84c510b6
193b6c49
d1526372
bfaeb554
b91029b8
7d499bdc
2b147f4b
fc75fb97
f50fc6c8
73979a33
1bde4038
29d4a60c
1445509a
46a8f581
66a8ea88
3344466a
6c9bea44
878b9dd6
144ef328
0c21d553
a7252cfd
0ab4fcd2
a4143713
f3f47340
ea5abdc7
eae7ce81
f4e605a4
76547fca
80c2e897
9e0b0f88
819479db
468b5b1c
5faca268
08fcb82f
cfd1fd81
0ba33b26
99e3bc42
89af90a3
c3f328ae
25ea0f0c
4faf223b
4cc9aa1f
b0e53a98
13452623
44f1594e
bd392929
aaec3ac6
dc421c82
153a3ce3
b698c156
c84c3143
500f23d4
fa00ffde
0d90efbf
5a9b4fb8
b89d09e8
5df6d5e4
38c0dcdb
c1a0a892
5fa7d197
b6a73613
c1d60c6b
44c25e0c
3bcc876f
b9d21f4e
e2c4572d
bf36e394
adc14bd5
74ade64b
39ecb177
de92b67d
2323205b
9aaddce5
21c67357
60e20c54
a203c51d
fa510f47
a02551dc
8caa24f6
68cab491
86d65427
466e54a8
088672bc
3048864c
85684807
628a7408
563d8f4a
abd65c1b
4f86c45f
7eec3ad6
130ecb62
2c6de871
50f9e314
111dcbe4
a25a85ac
5893e292
b38a6ece
c7632839
3dd3c04a
c6431ac3
59ce4068
b5032752
ba956719
76328603
0e0be5cc
c3686833
0e5de6a1
27fd9470
c6547183
a991c982
60753943
6e9565b0
1cb513c1
343aed9a
f490d13d
8e0f6f30
c63c928e
852728ad
5b1adc6b
e7a3d48d
1c4e3be0
4a15cdeb
1a779771
ef0ba5e9
709e9976
78baaea5
14ef1103
31f26bf4
eb7346b5
09423b27
1f8a2522
81515593
46a887ea
043a61b7
74745e2c
d342097c
119b1672
a118358c
c1a03742
03e59088
e28a7c68
9e44662a
25541fae
105862d7
78288f66
03400d3b
950ba323
3947721f
d1c14163
1d75acf1
44689149
93f00429
98e8886e
16113b90
d9245b69
371944ba
29f9acb8
99950d65
21152ab5
9f485fe4
e23d5910
a928e30a
3d5bdce0
9f8c6206
8952212b
02047772
dab1a0ac
777c5d8e
30eca8dc
ce8e4f0f
c11be311
f4b16ca3
ece700ff
2e630923
2dc673cf
2d4c7dd3
785ad2d8
e935c283
822026ae
60684a28
1c9dd491
55549136
4d4b64bb
64c68760
bc52276c
43b4e4f4
3e382f2a
6f04d33c
1d7aa314
817c2887
2a8b3a84
f5906889
b5a4d199
e2ecf30b
a3a06bd3
a27e4874
05ea2b35
fc6505b2
28c718da
110fa3a1
b9a09988
69149fa0
947cb08a
34167969
cfbe9472
2b97213a
e6c86435
159265c4
bdb253a3
ff080a0a
000000d9
00000000
04006fbc
04007024
0400708c
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000001
00000000
abcd330e
e66d1234
0005deec
0000000b
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000043
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00011b74
0000be18
00000000
0001fb1c
0002095c
0002070c
0002070c
0002070c
0002070c
0002070c
0002070c
0002070c
0002070c
0002070c
ffffffff
ffffffff
ffffffff
0000ffff
53410001
00494943
00000000
00000000
00000000
00000000
00000000
00000000
53410000
00494943
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
04007264
04007264
0400726c
0400726c
04007274
04007274
0400727c
0400727c
04007284
04007284
0400728c
0400728c
04007294
04007294
0400729c
0400729c
040072a4
040072a4
040072ac
040072ac
040072b4
040072b4
040072bc
040072bc
040072c4
040072c4
040072cc
040072cc
040072d4
040072d4
040072dc
040072dc
040072e4
040072e4
040072ec
040072ec
040072f4
040072f4
040072fc
040072fc
04007304
04007304
0400730c
0400730c
04007314
04007314
0400731c
0400731c
04007324
04007324
0400732c
0400732c
04007334
04007334
0400733c
0400733c
04007344
04007344
0400734c
0400734c
04007354
04007354
0400735c
0400735c
04007364
04007364
0400736c
0400736c
04007374
04007374
0400737c
0400737c
04007384
04007384
0400738c
0400738c
04007394
04007394
0400739c
0400739c
040073a4
040073a4
040073ac
040073ac
040073b4
040073b4
040073bc
040073bc
040073c4
040073c4
040073cc
040073cc
040073d4
040073d4
040073dc
040073dc
040073e4
040073e4
040073ec
040073ec
040073f4
040073f4
040073fc
040073fc
04007404
04007404
0400740c
0400740c
04007414
04007414
0400741c
0400741c
04007424
04007424
0400742c
0400742c
04007434
04007434
0400743c
0400743c
04007444
04007444
0400744c
0400744c
04007454
04007454
0400745c
0400745c
04007464
04007464
0400746c
0400746c
04007474
04007474
0400747c
0400747c
04007484
04007484
0400748c
0400748c
04007494
04007494
0400749c
0400749c
040074a4
040074a4
040074ac
040074ac
040074b4
040074b4
040074bc
040074bc
040074c4
040074c4
040074cc
040074cc
040074d4
040074d4
040074dc
040074dc
040074e4
040074e4
040074ec
040074ec
040074f4
040074f4
040074fc
040074fc
04007504
04007504
0400750c
0400750c
04007514
04007514
0400751c
0400751c
04007524
04007524
0400752c
0400752c
04007534
04007534
0400753c
0400753c
04007544
04007544
0400754c
0400754c
04007554
04007554
0400755c
0400755c
04007564
04007564
0400756c
0400756c
04007574
04007574
0400757c
0400757c
04007584
04007584
0400758c
0400758c
04007594
04007594
0400759c
0400759c
040075a4
040075a4
040075ac
040075ac
040075b4
040075b4
040075bc
040075bc
040075c4
040075c4
040075cc
040075cc
040075d4
040075d4
040075dc
040075dc
040075e4
040075e4
040075ec
040075ec
040075f4
040075f4
040075fc
040075fc
04007604
04007604
0400760c
0400760c
04007614
04007614
0400761c
0400761c
04007624
04007624
0400762c
0400762c
04007634
04007634
0400763c
0400763c
04007644
04007644
0400764c
0400764c
04007654
04007654
0400765c
0400765c
00000000
000207a0
04006cd0
ffffffff
00020000
00000010
00000000
00527a03
01017c01
00020d1b
00000048
00000018
fc00caec
000005c0
300e4400
8105936c
89028801
94049203
96079506
98099708
030b990a
c10a0254
c944c844
d444d344
d644d544
d844d744
d24cd944
44000e44
0000000b
0000004c
00000064
fc00d060
000004d0
300e4400
89028870
92018103
94059304
96079506
98099708
9a0b990a
010c030c
c844c10a
d244c944
d444d344
d644d544
d844d744
da44d944
44000e44
0000000b
00000000
10080100
0a030209
19201811
05040b12
211a130c
22293028
060d141b
1c150e07
38312a23
242b3239
170f161d
332c251e
2d343b3a
2e271f26
363d3c35
3f3e372f
00002a5c
00002b3c
00002a6c
00002b3c
00002b48
00002b3c
00002a6c
00002a5c
00002a5c
00002b48
00002a6c
00002a34
00002a34
00002a34
00002a74
02020100
03030303
04040404
04040404
05050505
05050505
05050505
05050505
06060606
06060606
06060606
06060606
06060606
06060606
06060606
06060606
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
20202000
20202020
28282020
20282828
20202020
20202020
20202020
20202020
10108820
10101010
10101010
10101010
04040410
04040404
10040404
10101010
41411010
41414141
01010101
01010101
01010101
01010101
01010101
10101010
42421010
42424242
02020202
02020202
02020202
02020202
02020202
10101010
00000020
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00005204
00004a40
00004a40
000051f8
00004a40
00004a40
00004a40
00004c2c
00004a40
00004a40
00005070
00005198
00004a40
00005088
000051b4
00004a40
000051a8
00004a10
00004a10
00004a10
00004a10
00004a10
00004a10
00004a10
00004a10
00004a10
00004a40
00004a40
00004a40
00004a40
00004a40
00004a40
00004a40
00004ca4
00004a40
00004fc8
00005294
00004ca4
00004ca4
00004ca4
00004a40
00004a40
00004a40
00004a40
00005288
00004a40
00004a40
0000521c
00004a40
00004a40
00004a40
00004ff0
00004a40
00005254
00004a40
00004a40
00005c64
00004a40
00004a40
00004a40
00004a40
00004a40
00004a40
00004a40
00004a40
00004ca4
00004a40
00004fc8
00005b24
00004ca4
00004ca4
00004ca4
00005184
00005b24
00004c6c
00004a40
000050dc
00004a40
00005094
00005c78
000050f0
00004c6c
00004a40
00004ff0
00004c64
00005bf8
00004a40
00004a40
00005c04
00004a40
00004c64
00006a6c
00006394
00006394
00006394
00006a54
00006a60
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006394
00006a54
00006a60
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
3fff8000
4a926576
153f804a
979ac94c
52028a20
7525c460
ce526a32
28ce329a
5de4a74d
3b5dc53d
5a929e8b
50ce526c
3d28f18b
0c17650d
75868175
4d48c976
58f89c66
5c54bc50
91c6cc65
a0aea60e
46a3e319
eab7851e
901b98fe
de8dddbb
ebfb9df9
4351aa7e
01370235
336c36b1
8cdfc66f
47c980e9
41a893ba
25fb50f8
6b71c76b
a6d53cbf
1f49ffcf
40d3c278
00000000
00000000
b59df020
ada82b70
40699dc5
00000000
00000000
00000000
c9bf0400
40348e1b
00000000
00000000
00000000
20000000
4019bebc
00000000
00000000
00000000
00000000
400c9c40
00000000
00000000
00000000
00000000
4005c800
00000000
00000000
00000000
00000000
4002a000
cffc2030
8123a1c3
9fde2de3
04c8d2ce
0ad8a6dd
d2cb8264
12d4f2ea
2de44925
534f3436
256bceae
f698f53f
01586bd3
c0bd87a6
82a5da57
32b5a2a6
04d4e731
d332e3f2
d21c7132
ee32db23
395a9049
5308a23e
1155fefb
1939fa91
4325637a
3cacc031
dbdee26d
b3f6d05d
e4a0ac7c
467c64bc
3e55ddd0
62242a20
98d747b3
e9a53f23
ea27a539
3f2aa87f
4af20b5b
18eda581
94ba67de
1ead4539
3f94cfb1
a9b3bf71
be687989
e15b4c2e
94bec44d
3fc9e695
7c3d3d4d
0d2b36ba
cefcfdc2
77118461
3fe4abcc
a4a8c155
6113404e
652bd3c3
1758e219
3ff1d1b7
70a3d70a
a3d70a3d
d70a3d70
0a3d70a3
3ff8a3d7
cccccccd
cccccccc
cccccccc
cccccccc
3ffbcccc
fffeffff
fff8fffc
ffe0fff0
ff80ffc0
fe00ff00
f800fc00
e000f000
8000c000
00000000
00000005
00000019
0000007d
00000000
00000000
3ff00000
00000000
40240000
00000000
40590000
00000000
408f4000
00000000
40c38800
00000000
40f86a00
00000000
412e8480
00000000
416312d0
00000000
4197d784
00000000
41cdcd65
20000000
4202a05f
e8000000
42374876
a2000000
426d1a94
e5400000
42a2309c
1e900000
42d6bcc4
26340000
430c6bf5
37e08000
4341c379
85d8a000
43763457
674ec800
43abc16d
60913d00
43e158e4
78b58c40
4415af1d
d6e2ef50
444b1ae4
064dd592
4480f0cf
c7e14af6
44b52d02
79d99db4
44ea7843
97d889bc
3c9cd2b2
d5a8a733
3949f623
44f4a73d
32a50ffd
cf8c979d
255bba08
64ac6f43
0ac80628
37e08000
4341c379
b5056e17
4693b8b5
e93ff9f5
4d384f03
f9301d32
5a827748
7f73bf3c
75154fdd
0000e90c
0000e178
0000e178
0000e900
0000e178
0000e178
0000e178
0000e31c
0000e178
0000e178
0000e758
0000e974
0000e178
0000e770
0000e930
0000e178
0000e924
0000e148
0000e148
0000e148
0000e148
0000e148
0000e148
0000e148
0000e148
0000e148
0000e178
0000e178
0000e178
0000e178
0000e178
0000e178
0000e178
0000e398
0000e178
0000e730
0000e984
0000e398
0000e398
0000e398
0000e178
0000e178
0000e178
0000e178
0000e8f4
0000e178
0000e178
0000e874
0000e178
0000e178
0000e178
0000e6b0
0000e178
0000e8c0
0000e178
0000e178
0000f3e0
0000e178
0000e178
0000e178
0000e178
0000e178
0000e178
0000e178
0000e178
0000e398
0000e178
0000e730
0000f278
0000e398
0000e398
0000e398
0000e8ac
0000f278
0000e360
0000e178
0000e7cc
0000e178
0000e77c
0000f3f4
0000e7e0
0000e360
0000e178
0000e6b0
0000e358
0000f334
0000e178
0000e178
0000f340
0000e178
0000e358
0000fdfc
0000fb40
0000fb40
0000fb40
0000fde4
0000fdf0
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fb40
0000fde4
0000fdf0
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
0001106c
00010ac0
00010ac0
00011060
00010ac0
00010ac0
00010ac0
00010c7c
00010ac0
00010ac0
00010fd8
000110d0
00010ac0
00010ffc
00011090
00010ac0
00011084
00010a88
00010a88
00010a88
00010a88
00010a88
00010a88
00010a88
00010a88
00010a88
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010f84
00010ccc
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010dc4
00010ac0
00010ac0
00010ac0
00010f44
00010ac0
00011030
00010ac0
00010ac0
0001187c
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010ac0
00010f84
00010cd0
00010ac0
00010ac0
00010ac0
0001101c
00010cd0
00010cc0
00010ac0
00011008
00010ac0
00011118
00010dc8
000110e0
00010cc0
00010ac0
00010f44
00010cb8
00011818
00010ac0
00010ac0
00011820
00010ac0
00010cb8
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
00012e9c
000128ac
000128ac
00012e90
000128ac
000128ac
000128ac
00012a18
000128ac
000128ac
00012e70
00012e60
000128ac
00012a7c
00012e20
000128ac
00012cb4
00012874
00012874
00012874
00012874
00012874
00012874
00012874
00012874
00012874
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
00012b50
00012d4c
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
00012d18
000128ac
000128ac
000128ac
00012afc
000128ac
00012ce8
000128ac
000128ac
00013590
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
000128ac
00012b50
00012b7c
000128ac
000128ac
000128ac
00012cd4
00012b7c
00012a60
000128ac
00012cc0
000128ac
00012c74
000135d8
00012c00
00012a60
000128ac
00012afc
00012a58
00013528
000128ac
000128ac
00013530
000128ac
00012a58
20202020
20202020
20202020
20202020
30303030
30303030
30303030
30303030
6f636544
676e6964
3a666f20
0a732520
00000000
4f525245
64203a52
646f6365
20676e69
6c696166
00006465
70616c45
20646573
656d6974
6625203a
00000a73
706d6f43
64657475
43504920
6625203a
0000000a
20555043
63746546
2e2e3a68
6625202e
000a2525
20555043
63657845
3a657475
6625202e
000a2525
20555043
6f6d654d
2e3a7972
6625202e
000a2525
78383025
0000203a
78323025
00000020
00206325
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
4952200a
562d4353
45504a20
65442047
69646f63
6220676e
68636e65
6b72616d
2b2b0a20
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
2b2b2b2b
000a2b2b
2067706a
78303233
20303432
00006b34
2067706a
78303233
20303432
00006b38
2067706a
78303233
20303432
006b3631
4f525245
49203a52
6c61766e
71206469
746e6175
74617a69
206e6f69
6c626174
44492065
6425203a
00000000
4f525245
49203a52
6c61766e
70206469
69636572
6e6f6973
00000000
00464e49
00666e69
004e414e
006e616e
33323130
37363534
62613938
66656463
00000000
33323130
37363534
42413938
46454443
00000000
6c756e28
0000296c
00000030
6e492d20
696e6966
00207974
666e4920
74696e69
00002079
004e614e
00642545
6c6c6142
7320636f
65636375
64656465
00000000
6d6f682f
62752f65
75746e75
636f442f
6e656d75
722f7374
76637369
756e672d
6f6f742d
6168636c
722f6e69
76637369
77656e2d
2f62696c
6c77656e
6c2f6269
2f636269
6c647473
6c2f6269
616f7464
0000632e
4e614e20
00000020
00000043
49534f50
00000058
0000002e
6d6f682f
62752f65
75746e75
636f442f
6e656d75
722f7374
76637369
756e672d
6f6f742d
6168636c
722f6e69
76637369
77656e2d
2f62696c
6c77656e
6c2f6269
2f636269
6c647473
6d2f6269
63657270
0000632e
7566202c
6974636e
203a6e6f
00000000
65737361
6f697472
2522206e
66202273
656c6961
66203a64
20656c69
22732522
696c202c
2520656e
25732564
00000a73
3dc7c5c4
3e43ef15
3e8e39da
3eb504f3
3ed4db31
3eec835e
3efb14be
3eb504f3
40273d74
3f8a8bd4
3f43ef15
3fb504f3
3fb504f3
3fec835e
04006cd0
00000000
4187d784
00000000
40590000
3eb504f3
3eec835e
3e43ef15
3e8e39da
3efb14be
3dc7c5c4
3ed4db31
3f43ef15
3fb504f3
40273d74
3f8a8bd4
3fb374bc
43000000
3eb020c5
3f36c8b4
3fe2d0e5
00000000
3ff00000
00000000
40240000
00000000
43500000
00000110
00018254
000000c8
